netcdf restart_out {
dimensions:
	mland = 1 ;
	mp_patch = 1 ;
	soil = 6 ;
	snow = 3 ;
	rad = 3 ;
	soil_carbon_pools = 2 ;
	plant_carbon_pools = 3 ;
	time = 1 ;
variables:
	double time(time) ;
		time:units = "seconds since 2002-01-01 00:00:00" ;
		time:coordinate = "LOC" ;
	float latitude(mland) ;
		latitude:units = "degrees_north" ;
	float longitude(mland) ;
		longitude:units = "degrees_east" ;
	float nap(mland) ;
		nap:long_name = "Number of active patches" ;
	float patchfrac(mp_patch) ;
		patchfrac:long_name = "Fraction of vegetated grid cell area occupied by a vegetation/soil patch" ;
	int mvtype ;
		mvtype:long_name = "Number of vegetation types" ;
	int mstype ;
		mstype:long_name = "Number of soil types" ;
	float tgg(soil, mp_patch) ;
		tgg:units = "K" ;
		tgg:long_name = "Average layer soil temperature" ;
		tgg:_FillValue = -1.e+33f ;
		tgg:missing_value = -1.e+33f ;
	double wb(soil, mp_patch) ;
		wb:units = "vol/vol" ;
		wb:long_name = "Average layer volumetric soil moisture" ;
		wb:_FillValue = -9.99999994495727e+32 ;
		wb:missing_value = -9.99999994495727e+32 ;
	double wbice(soil, mp_patch) ;
		wbice:units = "vol/vol" ;
		wbice:long_name = "Average layer volumetric soil ice" ;
		wbice:_FillValue = -9.99999994495727e+32 ;
		wbice:missing_value = -9.99999994495727e+32 ;
	float tss(mp_patch) ;
		tss:units = "K" ;
		tss:long_name = "Combined soil/snow temperature" ;
		tss:_FillValue = -1.e+33f ;
		tss:missing_value = -1.e+33f ;
	float albsoilsn(rad, mp_patch) ;
		albsoilsn:units = "-" ;
		albsoilsn:long_name = "Combined soil/snow albedo" ;
		albsoilsn:_FillValue = -1.e+33f ;
		albsoilsn:missing_value = -1.e+33f ;
	float rtsoil(mp_patch) ;
		rtsoil:units = "??" ;
		rtsoil:long_name = "Turbulent resistance for soil" ;
		rtsoil:_FillValue = -1.e+33f ;
		rtsoil:missing_value = -1.e+33f ;
	double gammzz(soil, mp_patch) ;
		gammzz:units = "J/kg/C" ;
		gammzz:long_name = "Heat capacity for each soil layer" ;
		gammzz:_FillValue = -9.99999994495727e+32 ;
		gammzz:missing_value = -9.99999994495727e+32 ;
	float runoff(mp_patch) ;
		runoff:units = "mm/timestep" ;
		runoff:long_name = "Total runoff" ;
		runoff:_FillValue = -1.e+33f ;
		runoff:missing_value = -1.e+33f ;
	float rnof1(mp_patch) ;
		rnof1:units = "mm/timestep" ;
		rnof1:long_name = "Surface runoff" ;
		rnof1:_FillValue = -1.e+33f ;
		rnof1:missing_value = -1.e+33f ;
	float rnof2(mp_patch) ;
		rnof2:units = "mm/timestep" ;
		rnof2:long_name = "Subsurface runoff" ;
		rnof2:_FillValue = -1.e+33f ;
		rnof2:missing_value = -1.e+33f ;
	float tggsn(snow, mp_patch) ;
		tggsn:units = "K" ;
		tggsn:long_name = "Average layer snow temperature" ;
		tggsn:_FillValue = -1.e+33f ;
		tggsn:missing_value = -1.e+33f ;
	float ssdnn(mp_patch) ;
		ssdnn:units = "kg/m^3" ;
		ssdnn:long_name = "Average snow density" ;
		ssdnn:_FillValue = -1.e+33f ;
		ssdnn:missing_value = -1.e+33f ;
	float ssdn(snow, mp_patch) ;
		ssdn:units = "kg/m^3" ;
		ssdn:long_name = "Average layer snow density" ;
		ssdn:_FillValue = -1.e+33f ;
		ssdn:missing_value = -1.e+33f ;
	float snowd(mp_patch) ;
		snowd:units = "mm" ;
		snowd:long_name = "Liquid water eqivalent snow depth" ;
		snowd:_FillValue = -1.e+33f ;
		snowd:missing_value = -1.e+33f ;
	float snage(mp_patch) ;
		snage:units = "??" ;
		snage:long_name = "Snow age" ;
		snage:_FillValue = -1.e+33f ;
		snage:missing_value = -1.e+33f ;
	float smass(snow, mp_patch) ;
		smass:units = "kg/m^2" ;
		smass:long_name = "Average layer snow mass" ;
		smass:_FillValue = -1.e+33f ;
		smass:missing_value = -1.e+33f ;
	float sdepth(snow, mp_patch) ;
		sdepth:units = "m" ;
		sdepth:long_name = "Snow layer depth" ;
		sdepth:_FillValue = -1.e+33f ;
		sdepth:missing_value = -1.e+33f ;
	float osnowd(mp_patch) ;
		osnowd:units = "mm" ;
		osnowd:long_name = "Previous time step snow depth in water equivalent" ;
		osnowd:_FillValue = -1.e+33f ;
		osnowd:missing_value = -1.e+33f ;
	int isflag(mp_patch) ;
		isflag:units = "-" ;
		isflag:long_name = "Snow layer scheme flag" ;
		isflag:_FillValue = -9999999 ;
		isflag:missing_value = -9999999 ;
	float cansto(mp_patch) ;
		cansto:units = "mm" ;
		cansto:long_name = "Canopy surface water storage" ;
		cansto:_FillValue = -1.e+33f ;
		cansto:missing_value = -1.e+33f ;
	float ghflux(mp_patch) ;
		ghflux:units = "W/m^2?" ;
		ghflux:long_name = "????" ;
		ghflux:_FillValue = -1.e+33f ;
		ghflux:missing_value = -1.e+33f ;
	float sghflux(mp_patch) ;
		sghflux:units = "W/m^2?" ;
		sghflux:long_name = "????" ;
		sghflux:_FillValue = -1.e+33f ;
		sghflux:missing_value = -1.e+33f ;
	float ga(mp_patch) ;
		ga:units = "W/m^2" ;
		ga:long_name = "Ground heat flux" ;
		ga:_FillValue = -1.e+33f ;
		ga:missing_value = -1.e+33f ;
	double dgdtg(mp_patch) ;
		dgdtg:units = "W/m^2/K" ;
		dgdtg:long_name = "Derivative of ground heat flux wrt soil temperature" ;
		dgdtg:_FillValue = -9.99999994495727e+32 ;
		dgdtg:missing_value = -9.99999994495727e+32 ;
	float fev(mp_patch) ;
		fev:units = "W/m^2" ;
		fev:long_name = "Latent heat flux from vegetation" ;
		fev:_FillValue = -1.e+33f ;
		fev:missing_value = -1.e+33f ;
	float fes(mp_patch) ;
		fes:units = "W/m^2" ;
		fes:long_name = "Latent heat flux from soil" ;
		fes:_FillValue = -1.e+33f ;
		fes:missing_value = -1.e+33f ;
	float fhs(mp_patch) ;
		fhs:units = "W/m^2" ;
		fhs:long_name = "Sensible heat flux from soil" ;
		fhs:_FillValue = -1.e+33f ;
		fhs:missing_value = -1.e+33f ;
	float cplant(plant_carbon_pools, mp_patch) ;
		cplant:units = "gC/m^2" ;
		cplant:long_name = "Plant carbon stores" ;
		cplant:_FillValue = -1.e+33f ;
		cplant:missing_value = -1.e+33f ;
	float csoil(soil_carbon_pools, mp_patch) ;
		csoil:units = "gC/m^2" ;
		csoil:long_name = "Soil carbon stores" ;
		csoil:_FillValue = -1.e+33f ;
		csoil:missing_value = -1.e+33f ;
	float wbtot0(mp_patch) ;
		wbtot0:units = "mm" ;
		wbtot0:long_name = "Initial time step soil water total" ;
		wbtot0:_FillValue = -1.e+33f ;
		wbtot0:missing_value = -1.e+33f ;
	float osnowd0(mp_patch) ;
		osnowd0:units = "mm" ;
		osnowd0:long_name = "Initial time step snow water total" ;
		osnowd0:_FillValue = -1.e+33f ;
		osnowd0:missing_value = -1.e+33f ;
	float albedo(rad, mp_patch) ;
		albedo:units = "-" ;
		albedo:long_name = "Albedo for shortwave and NIR radiation" ;
		albedo:_FillValue = -1.e+33f ;
		albedo:missing_value = -1.e+33f ;
	float trad(mp_patch) ;
		trad:units = "K" ;
		trad:long_name = "Surface radiative temperature (soil/snow/veg inclusive)" ;
		trad:_FillValue = -1.e+33f ;
		trad:missing_value = -1.e+33f ;
	int iveg(mp_patch) ;
		iveg:units = "-" ;
		iveg:long_name = "Vegetation type" ;
		iveg:_FillValue = -9999999 ;
		iveg:missing_value = -9999999 ;
	int isoil(mp_patch) ;
		isoil:units = "-" ;
		isoil:long_name = "Soil type" ;
		isoil:_FillValue = -9999999 ;
		isoil:missing_value = -9999999 ;
	float clay(mp_patch) ;
		clay:units = "-" ;
		clay:long_name = "Fraction of soil which is clay" ;
		clay:_FillValue = -1.e+33f ;
		clay:missing_value = -1.e+33f ;
	float sand(mp_patch) ;
		sand:units = "-" ;
		sand:long_name = "Fraction of soil which is sand" ;
		sand:_FillValue = -1.e+33f ;
		sand:missing_value = -1.e+33f ;
	float silt(mp_patch) ;
		silt:units = "-" ;
		silt:long_name = "Fraction of soil which is silt" ;
		silt:_FillValue = -1.e+33f ;
		silt:missing_value = -1.e+33f ;
	float ssat(mp_patch) ;
		ssat:units = "-" ;
		ssat:long_name = "Fraction of soil volume which is water @ saturation" ;
		ssat:_FillValue = -1.e+33f ;
		ssat:missing_value = -1.e+33f ;
	float sfc(mp_patch) ;
		sfc:units = "-" ;
		sfc:long_name = "Fraction of soil volume which is water @ field capacity" ;
		sfc:_FillValue = -1.e+33f ;
		sfc:missing_value = -1.e+33f ;
	float swilt(mp_patch) ;
		swilt:units = "-" ;
		swilt:long_name = "Fraction of soil volume which is water @ wilting point" ;
		swilt:_FillValue = -1.e+33f ;
		swilt:missing_value = -1.e+33f ;
	float zse(soil) ;
		zse:long_name = "Depth of each soil layer" ;
		zse:units = "m" ;
	float froot(soil, mp_patch) ;
		froot:units = "-" ;
		froot:long_name = "Fraction of roots in each soil layer" ;
		froot:_FillValue = -1.e+33f ;
		froot:missing_value = -1.e+33f ;
	float bch(mp_patch) ;
		bch:units = "-" ;
		bch:long_name = "Parameter b, Campbell eqn 1985" ;
		bch:_FillValue = -1.e+33f ;
		bch:missing_value = -1.e+33f ;
	float hyds(mp_patch) ;
		hyds:units = "m/s" ;
		hyds:long_name = "Hydraulic conductivity @ saturation" ;
		hyds:_FillValue = -1.e+33f ;
		hyds:missing_value = -1.e+33f ;
	float sucs(mp_patch) ;
		sucs:units = "m" ;
		sucs:long_name = "Suction @ saturation" ;
		sucs:_FillValue = -1.e+33f ;
		sucs:missing_value = -1.e+33f ;
	float css(mp_patch) ;
		css:units = "J/kg/C" ;
		css:long_name = "Heat capacity of soil minerals" ;
		css:_FillValue = -1.e+33f ;
		css:missing_value = -1.e+33f ;
	float rhosoil(mp_patch) ;
		rhosoil:units = "kg/m^3" ;
		rhosoil:long_name = "Density of soil minerals" ;
		rhosoil:_FillValue = -1.e+33f ;
		rhosoil:missing_value = -1.e+33f ;
	float rs20(mp_patch) ;
		rs20:units = "-" ;
		rs20:long_name = "Soil respiration coefficient at 20C" ;
		rs20:_FillValue = -1.e+33f ;
		rs20:missing_value = -1.e+33f ;
	float albsoil(rad, mp_patch) ;
		albsoil:units = "-" ;
		albsoil:long_name = "Soil reflectance" ;
		albsoil:_FillValue = -1.e+33f ;
		albsoil:missing_value = -1.e+33f ;
	float hc(mp_patch) ;
		hc:units = "m" ;
		hc:long_name = "Height of canopy" ;
		hc:_FillValue = -1.e+33f ;
		hc:missing_value = -1.e+33f ;
	float canst1(mp_patch) ;
		canst1:units = "mm/LAI" ;
		canst1:long_name = "Max water intercepted by canopy" ;
		canst1:_FillValue = -1.e+33f ;
		canst1:missing_value = -1.e+33f ;
	float dleaf(mp_patch) ;
		dleaf:units = "m" ;
		dleaf:long_name = "Chararacteristic length of leaf" ;
		dleaf:_FillValue = -1.e+33f ;
		dleaf:missing_value = -1.e+33f ;
	float frac4(mp_patch) ;
		frac4:units = "-" ;
		frac4:long_name = "Fraction of plants which are C4" ;
		frac4:_FillValue = -1.e+33f ;
		frac4:missing_value = -1.e+33f ;
	float ejmax(mp_patch) ;
		ejmax:units = "mol/m^2/s" ;
		ejmax:long_name = "Max potential electron transport rate top leaf" ;
		ejmax:_FillValue = -1.e+33f ;
		ejmax:missing_value = -1.e+33f ;
	float vcmax(mp_patch) ;
		vcmax:units = "mol/m^2/s" ;
		vcmax:long_name = "Maximum RuBP carboxylation rate top leaf" ;
		vcmax:_FillValue = -1.e+33f ;
		vcmax:missing_value = -1.e+33f ;
	float rp20(mp_patch) ;
		rp20:units = "-" ;
		rp20:long_name = "Plant respiration coefficient at 20C" ;
		rp20:_FillValue = -1.e+33f ;
		rp20:missing_value = -1.e+33f ;
	float rpcoef(mp_patch) ;
		rpcoef:units = "1/C" ;
		rpcoef:long_name = "Temperature coef nonleaf plant respiration" ;
		rpcoef:_FillValue = -1.e+33f ;
		rpcoef:missing_value = -1.e+33f ;
	float shelrb(mp_patch) ;
		shelrb:units = "-" ;
		shelrb:long_name = "Sheltering factor" ;
		shelrb:_FillValue = -1.e+33f ;
		shelrb:missing_value = -1.e+33f ;
	float xfang(mp_patch) ;
		xfang:units = "-" ;
		xfang:long_name = "Leaf angle parameter" ;
		xfang:_FillValue = -1.e+33f ;
		xfang:missing_value = -1.e+33f ;
	float wai(mp_patch) ;
		wai:units = "-" ;
		wai:long_name = "Wood area index" ;
		wai:_FillValue = -1.e+33f ;
		wai:missing_value = -1.e+33f ;
	float vegcf(mp_patch) ;
		vegcf:units = "-" ;
		vegcf:long_name = "vegcf" ;
		vegcf:_FillValue = -1.e+33f ;
		vegcf:missing_value = -1.e+33f ;
	float extkn(mp_patch) ;
		extkn:units = "-" ;
		extkn:long_name = "Extinction coef for vertical nitrogen profile" ;
		extkn:_FillValue = -1.e+33f ;
		extkn:missing_value = -1.e+33f ;
	float tminvj(mp_patch) ;
		tminvj:units = "C" ;
		tminvj:long_name = "Min temperature for the start of photosynthesis" ;
		tminvj:_FillValue = -1.e+33f ;
		tminvj:missing_value = -1.e+33f ;
	float tmaxvj(mp_patch) ;
		tmaxvj:units = "C" ;
		tmaxvj:long_name = "Max temperature for the start of photosynthesis" ;
		tmaxvj:_FillValue = -1.e+33f ;
		tmaxvj:missing_value = -1.e+33f ;
	float vbeta(mp_patch) ;
		vbeta:units = "-" ;
		vbeta:long_name = "Stomatal sensitivity to soil water" ;
		vbeta:_FillValue = -1.e+33f ;
		vbeta:missing_value = -1.e+33f ;
	float xalbnir(mp_patch) ;
		xalbnir:units = "-" ;
		xalbnir:long_name = "modifier for albedo in near ir band" ;
		xalbnir:_FillValue = -1.e+33f ;
		xalbnir:missing_value = -1.e+33f ;
	float ratecp(plant_carbon_pools) ;
		ratecp:long_name = "Plant carbon rate constant" ;
		ratecp:units = "1/year" ;
	float ratecs(soil_carbon_pools) ;
		ratecs:long_name = "Soil carbon rate constant" ;
		ratecs:units = "1/year" ;
	int meth(mp_patch) ;
		meth:units = "-" ;
		meth:long_name = "Canopy turbulence parameterisation switch" ;
		meth:_FillValue = -9999999 ;
		meth:missing_value = -9999999 ;
	float za_uv(mp_patch) ;
		za_uv:units = "m" ;
		za_uv:long_name = "Reference height (lowest atm. model layer) for momentum" ;
		za_uv:_FillValue = -1.e+33f ;
		za_uv:missing_value = -1.e+33f ;
	float za_tq(mp_patch) ;
		za_tq:units = "m" ;
		za_tq:long_name = "Reference height (lowest atm. model layer) for scalars" ;
		za_tq:_FillValue = -1.e+33f ;
		za_tq:missing_value = -1.e+33f ;

// global attributes:
		:Production = "2012/12/19 at 01:33:42" ;
		:Source = "CABLE LSM restart file" ;
		:CABLE_input_file = "/projects/access/CABLE-AUX/offline/TumbaFluxnet.1.3_met.nc" ;
data:

 time = 126232200 ;

 latitude = -35.656 ;

 longitude = 148.15 ;

 nap = 1 ;

 patchfrac = 1 ;

 mvtype = 17 ;

 mstype = 9 ;

 tgg =
  297.3815,
  300.227,
  301.2762,
  293.7083,
  286.6244,
  282.3425 ;

 wb =
  0.0768643620487479,
  0.15367652072873,
  0.183915351659266,
  0.246320550657871,
  0.287873155154424,
  0.320297168821936 ;

 wbice =
  0,
  0,
  0,
  0,
  0,
  0 ;

 tss = 297.3815 ;

 albsoilsn =
  0.05869506,
  0.1173901,
  0 ;

 rtsoil = 67.80319 ;

 gammzz =
  28153.9938474447,
  80858.6067915507,
  234329.005582272,
  729990.739733053,
  2126800.49506748,
  6022452.49501962 ;

 runoff = 0.01260123 ;

 rnof1 = 0 ;

 rnof2 = 0.01260123 ;

 tggsn =
  273.16,
  273.16,
  273.16 ;

 ssdnn = 120 ;

 ssdn =
  120,
  120,
  120 ;

 snowd = 0 ;

 snage = 0 ;

 smass =
  0,
  0,
  0 ;

 sdepth =
  0,
  0,
  0 ;

 osnowd = 0 ;

 isflag = 0 ;

 cansto = 0 ;

 ghflux = -40.04517 ;

 sghflux = 0 ;

 ga = -123.5866 ;

 dgdtg = -21.4920120239258 ;

 fev = 13.9204 ;

 fes = 0.1569544 ;

 fhs = 70.47467 ;

 cplant =
  213.262,
  15272.16,
  1167.961 ;

 csoil =
  7650.634,
  1114.739 ;

 wbtot0 = 1077.444 ;

 osnowd0 = 0 ;

 albedo =
  0.02499556,
  0.114129,
  0 ;

 trad = 295.4286 ;

 iveg = 2 ;

 isoil = 2 ;

 clay = 0.3 ;

 sand = 0.37 ;

 silt = 0.33 ;

 ssat = 0.4171363 ;

 sfc = 0.2644416 ;

 swilt = 0.1536539 ;

 zse = 0.022, 0.058, 0.154, 0.409, 1.085, 2.872 ;

 froot =
  0.08169878,
  0.1848004,
  0.3295795,
  0.3210971,
  0.08158642,
  0.00123781 ;

 bch = 7.03 ;

 hyds = 5.984919e-06 ;

 sucs = -0.1365896 ;

 css = 813.1797 ;

 rhosoil = 1573.732 ;

 rs20 = 1 ;

 albsoil =
  0.08804259,
  0.1760852,
  0 ;

 hc = 45 ;

 canst1 = 0.1 ;

 dleaf = 0.07071068 ;

 frac4 = 0 ;

 ejmax = 0.00011 ;

 vcmax = 5.5e-05 ;

 rp20 = 0.6 ;

 rpcoef = 0.0832 ;

 shelrb = 2 ;

 xfang = 0.1 ;

 wai = 1 ;

 vegcf = 14 ;

 extkn = 0.001 ;

 tminvj = -15 ;

 tmaxvj = -10 ;

 vbeta = 2 ;

 xalbnir = 1 ;

 ratecp = 1, 0.03, 0.14 ;

 ratecs = 2, 0.5 ;

 meth = 1 ;

 za_uv = 70 ;

 za_tq = 70 ;
}
