netcdf Loobos_1997 {
dimensions:
	time = UNLIMITED ; // (17520 currently)
	z = 4 ;
	y = 1 ;
	x = 1 ;
variables:
	double iveg(z, y, x) ;
		iveg:units = "-" ;
		iveg:missing_value = -9999.f ;
		iveg:long_name = "Vegetation type" ;
	double patchfrac(z, y, x) ;
		patchfrac:units = "-" ;
		patchfrac:missing_value = -9999.f ;
		patchfrac:long_name = "Vegetation type" ;
	double time(time) ;
		time:units = "seconds since 1996-12-31 23:30:00" ;
		time:long_name = "time" ;
		time:calendar = "standard" ;
	double z(z) ;
		z:long_name = "z dimension" ;
	double y(y) ;
		y:long_name = "y dimension" ;
	double x(x) ;
		x:long_name = "x dimension" ;
	double latitude(y, x) ;
		latitude:units = "degrees_north" ;
		latitude:missing_value = -9999. ;
		latitude:long_name = "Latitude" ;
	double longitude(y, x) ;
		longitude:units = "degrees_east" ;
		longitude:missing_value = -9999. ;
		longitude:long_name = "Longitude" ;
	double SWdown(time, y, x) ;
		SWdown:units = "W/m^2" ;
		SWdown:missing_value = -9999. ;
		SWdown:long_name = "Surface incident shortwave radiation" ;
		SWdown:CF_name = "surface_downwelling_shortwave_flux_in_air" ;
	double Tair(time, z, y, x) ;
		Tair:units = "K" ;
		Tair:missing_value = -9999. ;
		Tair:long_name = "Near surface air temperature" ;
		Tair:CF_name = "surface_temperature" ;
	double Rainf(time, y, x) ;
		Rainf:units = "mm/s" ;
		Rainf:missing_value = -9999. ;
		Rainf:long_name = "Rainfall rate" ;
		Rainf:CF_name = "precipitation_flux" ;
	double Snowf(time, y, x) ;
		Snowf:units = "mm/s" ;
		Snowf:missing_value = -9999. ;
		Snowf:long_name = "Snowfall rate" ;
		Snowf:CF_name = "snowfall_flux" ;
	double Qair(time, z, y, x) ;
		Qair:units = "kg/kg" ;
		Qair:missing_value = -9999. ;
		Qair:long_name = "Near surface specific humidity" ;
		Qair:CF_name = "surface_specific_humidity" ;
	double Wind(time, z, y, x) ;
		Wind:units = "m/s" ;
		Wind:missing_value = -9999. ;
		Wind:long_name = "Scalar windspeed" ;
		Wind:CF_name = "wind_speed" ;
	double PSurf(time, y, x) ;
		PSurf:units = "Pa" ;
		PSurf:missing_value = -9999. ;
		PSurf:long_name = "Surface air pressure" ;
		PSurf:CF_name = "surface_air_pressure" ;
	double LWdown(time, y, x) ;
		LWdown:units = "W/m^2" ;
		LWdown:missing_value = -9999. ;
		LWdown:long_name = "Surface incident longwave radiation" ;
		LWdown:CF_name = "surface_downwelling_longwave_flux_in_air" ;
	double CO2air(time, z, y, x) ;
		CO2air:units = "ppm" ;
		CO2air:missing_value = -9999. ;
		CO2air:long_name = "" ;
		CO2air:CF_name = "" ;
	double hc(y, x) ;
		hc:units = "m" ;
		hc:missing_value = -9999. ;
		hc:long_name = "canopy height" ;
	double za(y, x) ;
		za:units = "m" ;
		za:missing_value = -9999. ;
		za:long_name = "reference height" ;

// global attributes:
		:description = "Loobos met data, created by Martin De Kauwe" ;
		:history = "Created by: generate_CABLE_netcdf_met.py" ;
		:creation_date = "2019-11-14 12:32:16.113395" ;
		:contact = "mdekauwe@gmail.com" ;
		:_NCProperties = "version=2,netcdf=4.7.0,hdf5=1.10.5" ;
data:

 iveg =
  1,
  2,
  6,
  14 ;

 patchfrac =
  0.355,
  0.355,
  0.208,
  0.082 ;

 time = 0, 1800, 3600, 5400, 7200, 9000, 10800, 12600, 14400, 16200, 18000, 
    19800, 21600, 23400, 25200, 27000, 28800, 30600, 32400, 34200, 36000, 
    37800, 39600, 41400, 43200, 45000, 46800, 48600, 50400, 52200, 54000, 
    55800, 57600, 59400, 61200, 63000, 64800, 66600, 68400, 70200, 72000, 
    73800, 75600, 77400, 79200, 81000, 82800, 84600, 86400, 88200, 90000, 
    91800, 93600, 95400, 97200, 99000, 100800, 102600, 104400, 106200, 
    108000, 109800, 111600, 113400, 115200, 117000, 118800, 120600, 122400, 
    124200, 126000, 127800, 129600, 131400, 133200, 135000, 136800, 138600, 
    140400, 142200, 144000, 145800, 147600, 149400, 151200, 153000, 154800, 
    156600, 158400, 160200, 162000, 163800, 165600, 167400, 169200, 171000, 
    172800, 174600, 176400, 178200, 180000, 181800, 183600, 185400, 187200, 
    189000, 190800, 192600, 194400, 196200, 198000, 199800, 201600, 203400, 
    205200, 207000, 208800, 210600, 212400, 214200, 216000, 217800, 219600, 
    221400, 223200, 225000, 226800, 228600, 230400, 232200, 234000, 235800, 
    237600, 239400, 241200, 243000, 244800, 246600, 248400, 250200, 252000, 
    253800, 255600, 257400, 259200, 261000, 262800, 264600, 266400, 268200, 
    270000, 271800, 273600, 275400, 277200, 279000, 280800, 282600, 284400, 
    286200, 288000, 289800, 291600, 293400, 295200, 297000, 298800, 300600, 
    302400, 304200, 306000, 307800, 309600, 311400, 313200, 315000, 316800, 
    318600, 320400, 322200, 324000, 325800, 327600, 329400, 331200, 333000, 
    334800, 336600, 338400, 340200, 342000, 343800, 345600, 347400, 349200, 
    351000, 352800, 354600, 356400, 358200, 360000, 361800, 363600, 365400, 
    367200, 369000, 370800, 372600, 374400, 376200, 378000, 379800, 381600, 
    383400, 385200, 387000, 388800, 390600, 392400, 394200, 396000, 397800, 
    399600, 401400, 403200, 405000, 406800, 408600, 410400, 412200, 414000, 
    415800, 417600, 419400, 421200, 423000, 424800, 426600, 428400, 430200, 
    432000, 433800, 435600, 437400, 439200, 441000, 442800, 444600, 446400, 
    448200, 450000, 451800, 453600, 455400, 457200, 459000, 460800, 462600, 
    464400, 466200, 468000, 469800, 471600, 473400, 475200, 477000, 478800, 
    480600, 482400, 484200, 486000, 487800, 489600, 491400, 493200, 495000, 
    496800, 498600, 500400, 502200, 504000, 505800, 507600, 509400, 511200, 
    513000, 514800, 516600, 518400, 520200, 522000, 523800, 525600, 527400, 
    529200, 531000, 532800, 534600, 536400, 538200, 540000, 541800, 543600, 
    545400, 547200, 549000, 550800, 552600, 554400, 556200, 558000, 559800, 
    561600, 563400, 565200, 567000, 568800, 570600, 572400, 574200, 576000, 
    577800, 579600, 581400, 583200, 585000, 586800, 588600, 590400, 592200, 
    594000, 595800, 597600, 599400, 601200, 603000, 604800, 606600, 608400, 
    610200, 612000, 613800, 615600, 617400, 619200, 621000, 622800, 624600, 
    626400, 628200, 630000, 631800, 633600, 635400, 637200, 639000, 640800, 
    642600, 644400, 646200, 648000, 649800, 651600, 653400, 655200, 657000, 
    658800, 660600, 662400, 664200, 666000, 667800, 669600, 671400, 673200, 
    675000, 676800, 678600, 680400, 682200, 684000, 685800, 687600, 689400, 
    691200, 693000, 694800, 696600, 698400, 700200, 702000, 703800, 705600, 
    707400, 709200, 711000, 712800, 714600, 716400, 718200, 720000, 721800, 
    723600, 725400, 727200, 729000, 730800, 732600, 734400, 736200, 738000, 
    739800, 741600, 743400, 745200, 747000, 748800, 750600, 752400, 754200, 
    756000, 757800, 759600, 761400, 763200, 765000, 766800, 768600, 770400, 
    772200, 774000, 775800, 777600, 779400, 781200, 783000, 784800, 786600, 
    788400, 790200, 792000, 793800, 795600, 797400, 799200, 801000, 802800, 
    804600, 806400, 808200, 810000, 811800, 813600, 815400, 817200, 819000, 
    820800, 822600, 824400, 826200, 828000, 829800, 831600, 833400, 835200, 
    837000, 838800, 840600, 842400, 844200, 846000, 847800, 849600, 851400, 
    853200, 855000, 856800, 858600, 860400, 862200, 864000, 865800, 867600, 
    869400, 871200, 873000, 874800, 876600, 878400, 880200, 882000, 883800, 
    885600, 887400, 889200, 891000, 892800, 894600, 896400, 898200, 900000, 
    901800, 903600, 905400, 907200, 909000, 910800, 912600, 914400, 916200, 
    918000, 919800, 921600, 923400, 925200, 927000, 928800, 930600, 932400, 
    934200, 936000, 937800, 939600, 941400, 943200, 945000, 946800, 948600, 
    950400, 952200, 954000, 955800, 957600, 959400, 961200, 963000, 964800, 
    966600, 968400, 970200, 972000, 973800, 975600, 977400, 979200, 981000, 
    982800, 984600, 986400, 988200, 990000, 991800, 993600, 995400, 997200, 
    999000, 1000800, 1002600, 1004400, 1006200, 1008000, 1009800, 1011600, 
    1013400, 1015200, 1017000, 1018800, 1020600, 1022400, 1024200, 1026000, 
    1027800, 1029600, 1031400, 1033200, 1035000, 1036800, 1038600, 1040400, 
    1042200, 1044000, 1045800, 1047600, 1049400, 1051200, 1053000, 1054800, 
    1056600, 1058400, 1060200, 1062000, 1063800, 1065600, 1067400, 1069200, 
    1071000, 1072800, 1074600, 1076400, 1078200, 1080000, 1081800, 1083600, 
    1085400, 1087200, 1089000, 1090800, 1092600, 1094400, 1096200, 1098000, 
    1099800, 1101600, 1103400, 1105200, 1107000, 1108800, 1110600, 1112400, 
    1114200, 1116000, 1117800, 1119600, 1121400, 1123200, 1125000, 1126800, 
    1128600, 1130400, 1132200, 1134000, 1135800, 1137600, 1139400, 1141200, 
    1143000, 1144800, 1146600, 1148400, 1150200, 1152000, 1153800, 1155600, 
    1157400, 1159200, 1161000, 1162800, 1164600, 1166400, 1168200, 1170000, 
    1171800, 1173600, 1175400, 1177200, 1179000, 1180800, 1182600, 1184400, 
    1186200, 1188000, 1189800, 1191600, 1193400, 1195200, 1197000, 1198800, 
    1200600, 1202400, 1204200, 1206000, 1207800, 1209600, 1211400, 1213200, 
    1215000, 1216800, 1218600, 1220400, 1222200, 1224000, 1225800, 1227600, 
    1229400, 1231200, 1233000, 1234800, 1236600, 1238400, 1240200, 1242000, 
    1243800, 1245600, 1247400, 1249200, 1251000, 1252800, 1254600, 1256400, 
    1258200, 1260000, 1261800, 1263600, 1265400, 1267200, 1269000, 1270800, 
    1272600, 1274400, 1276200, 1278000, 1279800, 1281600, 1283400, 1285200, 
    1287000, 1288800, 1290600, 1292400, 1294200, 1296000, 1297800, 1299600, 
    1301400, 1303200, 1305000, 1306800, 1308600, 1310400, 1312200, 1314000, 
    1315800, 1317600, 1319400, 1321200, 1323000, 1324800, 1326600, 1328400, 
    1330200, 1332000, 1333800, 1335600, 1337400, 1339200, 1341000, 1342800, 
    1344600, 1346400, 1348200, 1350000, 1351800, 1353600, 1355400, 1357200, 
    1359000, 1360800, 1362600, 1364400, 1366200, 1368000, 1369800, 1371600, 
    1373400, 1375200, 1377000, 1378800, 1380600, 1382400, 1384200, 1386000, 
    1387800, 1389600, 1391400, 1393200, 1395000, 1396800, 1398600, 1400400, 
    1402200, 1404000, 1405800, 1407600, 1409400, 1411200, 1413000, 1414800, 
    1416600, 1418400, 1420200, 1422000, 1423800, 1425600, 1427400, 1429200, 
    1431000, 1432800, 1434600, 1436400, 1438200, 1440000, 1441800, 1443600, 
    1445400, 1447200, 1449000, 1450800, 1452600, 1454400, 1456200, 1458000, 
    1459800, 1461600, 1463400, 1465200, 1467000, 1468800, 1470600, 1472400, 
    1474200, 1476000, 1477800, 1479600, 1481400, 1483200, 1485000, 1486800, 
    1488600, 1490400, 1492200, 1494000, 1495800, 1497600, 1499400, 1501200, 
    1503000, 1504800, 1506600, 1508400, 1510200, 1512000, 1513800, 1515600, 
    1517400, 1519200, 1521000, 1522800, 1524600, 1526400, 1528200, 1530000, 
    1531800, 1533600, 1535400, 1537200, 1539000, 1540800, 1542600, 1544400, 
    1546200, 1548000, 1549800, 1551600, 1553400, 1555200, 1557000, 1558800, 
    1560600, 1562400, 1564200, 1566000, 1567800, 1569600, 1571400, 1573200, 
    1575000, 1576800, 1578600, 1580400, 1582200, 1584000, 1585800, 1587600, 
    1589400, 1591200, 1593000, 1594800, 1596600, 1598400, 1600200, 1602000, 
    1603800, 1605600, 1607400, 1609200, 1611000, 1612800, 1614600, 1616400, 
    1618200, 1620000, 1621800, 1623600, 1625400, 1627200, 1629000, 1630800, 
    1632600, 1634400, 1636200, 1638000, 1639800, 1641600, 1643400, 1645200, 
    1647000, 1648800, 1650600, 1652400, 1654200, 1656000, 1657800, 1659600, 
    1661400, 1663200, 1665000, 1666800, 1668600, 1670400, 1672200, 1674000, 
    1675800, 1677600, 1679400, 1681200, 1683000, 1684800, 1686600, 1688400, 
    1690200, 1692000, 1693800, 1695600, 1697400, 1699200, 1701000, 1702800, 
    1704600, 1706400, 1708200, 1710000, 1711800, 1713600, 1715400, 1717200, 
    1719000, 1720800, 1722600, 1724400, 1726200, 1728000, 1729800, 1731600, 
    1733400, 1735200, 1737000, 1738800, 1740600, 1742400, 1744200, 1746000, 
    1747800, 1749600, 1751400, 1753200, 1755000, 1756800, 1758600, 1760400, 
    1762200, 1764000, 1765800, 1767600, 1769400, 1771200, 1773000, 1774800, 
    1776600, 1778400, 1780200, 1782000, 1783800, 1785600, 1787400, 1789200, 
    1791000, 1792800, 1794600, 1796400, 1798200, 1800000, 1801800, 1803600, 
    1805400, 1807200, 1809000, 1810800, 1812600, 1814400, 1816200, 1818000, 
    1819800, 1821600, 1823400, 1825200, 1827000, 1828800, 1830600, 1832400, 
    1834200, 1836000, 1837800, 1839600, 1841400, 1843200, 1845000, 1846800, 
    1848600, 1850400, 1852200, 1854000, 1855800, 1857600, 1859400, 1861200, 
    1863000, 1864800, 1866600, 1868400, 1870200, 1872000, 1873800, 1875600, 
    1877400, 1879200, 1881000, 1882800, 1884600, 1886400, 1888200, 1890000, 
    1891800, 1893600, 1895400, 1897200, 1899000, 1900800, 1902600, 1904400, 
    1906200, 1908000, 1909800, 1911600, 1913400, 1915200, 1917000, 1918800, 
    1920600, 1922400, 1924200, 1926000, 1927800, 1929600, 1931400, 1933200, 
    1935000, 1936800, 1938600, 1940400, 1942200, 1944000, 1945800, 1947600, 
    1949400, 1951200, 1953000, 1954800, 1956600, 1958400, 1960200, 1962000, 
    1963800, 1965600, 1967400, 1969200, 1971000, 1972800, 1974600, 1976400, 
    1978200, 1980000, 1981800, 1983600, 1985400, 1987200, 1989000, 1990800, 
    1992600, 1994400, 1996200, 1998000, 1999800, 2001600, 2003400, 2005200, 
    2007000, 2008800, 2010600, 2012400, 2014200, 2016000, 2017800, 2019600, 
    2021400, 2023200, 2025000, 2026800, 2028600, 2030400, 2032200, 2034000, 
    2035800, 2037600, 2039400, 2041200, 2043000, 2044800, 2046600, 2048400, 
    2050200, 2052000, 2053800, 2055600, 2057400, 2059200, 2061000, 2062800, 
    2064600, 2066400, 2068200, 2070000, 2071800, 2073600, 2075400, 2077200, 
    2079000, 2080800, 2082600, 2084400, 2086200, 2088000, 2089800, 2091600, 
    2093400, 2095200, 2097000, 2098800, 2100600, 2102400, 2104200, 2106000, 
    2107800, 2109600, 2111400, 2113200, 2115000, 2116800, 2118600, 2120400, 
    2122200, 2124000, 2125800, 2127600, 2129400, 2131200, 2133000, 2134800, 
    2136600, 2138400, 2140200, 2142000, 2143800, 2145600, 2147400, 2149200, 
    2151000, 2152800, 2154600, 2156400, 2158200, 2160000, 2161800, 2163600, 
    2165400, 2167200, 2169000, 2170800, 2172600, 2174400, 2176200, 2178000, 
    2179800, 2181600, 2183400, 2185200, 2187000, 2188800, 2190600, 2192400, 
    2194200, 2196000, 2197800, 2199600, 2201400, 2203200, 2205000, 2206800, 
    2208600, 2210400, 2212200, 2214000, 2215800, 2217600, 2219400, 2221200, 
    2223000, 2224800, 2226600, 2228400, 2230200, 2232000, 2233800, 2235600, 
    2237400, 2239200, 2241000, 2242800, 2244600, 2246400, 2248200, 2250000, 
    2251800, 2253600, 2255400, 2257200, 2259000, 2260800, 2262600, 2264400, 
    2266200, 2268000, 2269800, 2271600, 2273400, 2275200, 2277000, 2278800, 
    2280600, 2282400, 2284200, 2286000, 2287800, 2289600, 2291400, 2293200, 
    2295000, 2296800, 2298600, 2300400, 2302200, 2304000, 2305800, 2307600, 
    2309400, 2311200, 2313000, 2314800, 2316600, 2318400, 2320200, 2322000, 
    2323800, 2325600, 2327400, 2329200, 2331000, 2332800, 2334600, 2336400, 
    2338200, 2340000, 2341800, 2343600, 2345400, 2347200, 2349000, 2350800, 
    2352600, 2354400, 2356200, 2358000, 2359800, 2361600, 2363400, 2365200, 
    2367000, 2368800, 2370600, 2372400, 2374200, 2376000, 2377800, 2379600, 
    2381400, 2383200, 2385000, 2386800, 2388600, 2390400, 2392200, 2394000, 
    2395800, 2397600, 2399400, 2401200, 2403000, 2404800, 2406600, 2408400, 
    2410200, 2412000, 2413800, 2415600, 2417400, 2419200, 2421000, 2422800, 
    2424600, 2426400, 2428200, 2430000, 2431800, 2433600, 2435400, 2437200, 
    2439000, 2440800, 2442600, 2444400, 2446200, 2448000, 2449800, 2451600, 
    2453400, 2455200, 2457000, 2458800, 2460600, 2462400, 2464200, 2466000, 
    2467800, 2469600, 2471400, 2473200, 2475000, 2476800, 2478600, 2480400, 
    2482200, 2484000, 2485800, 2487600, 2489400, 2491200, 2493000, 2494800, 
    2496600, 2498400, 2500200, 2502000, 2503800, 2505600, 2507400, 2509200, 
    2511000, 2512800, 2514600, 2516400, 2518200, 2520000, 2521800, 2523600, 
    2525400, 2527200, 2529000, 2530800, 2532600, 2534400, 2536200, 2538000, 
    2539800, 2541600, 2543400, 2545200, 2547000, 2548800, 2550600, 2552400, 
    2554200, 2556000, 2557800, 2559600, 2561400, 2563200, 2565000, 2566800, 
    2568600, 2570400, 2572200, 2574000, 2575800, 2577600, 2579400, 2581200, 
    2583000, 2584800, 2586600, 2588400, 2590200, 2592000, 2593800, 2595600, 
    2597400, 2599200, 2601000, 2602800, 2604600, 2606400, 2608200, 2610000, 
    2611800, 2613600, 2615400, 2617200, 2619000, 2620800, 2622600, 2624400, 
    2626200, 2628000, 2629800, 2631600, 2633400, 2635200, 2637000, 2638800, 
    2640600, 2642400, 2644200, 2646000, 2647800, 2649600, 2651400, 2653200, 
    2655000, 2656800, 2658600, 2660400, 2662200, 2664000, 2665800, 2667600, 
    2669400, 2671200, 2673000, 2674800, 2676600, 2678400, 2680200, 2682000, 
    2683800, 2685600, 2687400, 2689200, 2691000, 2692800, 2694600, 2696400, 
    2698200, 2700000, 2701800, 2703600, 2705400, 2707200, 2709000, 2710800, 
    2712600, 2714400, 2716200, 2718000, 2719800, 2721600, 2723400, 2725200, 
    2727000, 2728800, 2730600, 2732400, 2734200, 2736000, 2737800, 2739600, 
    2741400, 2743200, 2745000, 2746800, 2748600, 2750400, 2752200, 2754000, 
    2755800, 2757600, 2759400, 2761200, 2763000, 2764800, 2766600, 2768400, 
    2770200, 2772000, 2773800, 2775600, 2777400, 2779200, 2781000, 2782800, 
    2784600, 2786400, 2788200, 2790000, 2791800, 2793600, 2795400, 2797200, 
    2799000, 2800800, 2802600, 2804400, 2806200, 2808000, 2809800, 2811600, 
    2813400, 2815200, 2817000, 2818800, 2820600, 2822400, 2824200, 2826000, 
    2827800, 2829600, 2831400, 2833200, 2835000, 2836800, 2838600, 2840400, 
    2842200, 2844000, 2845800, 2847600, 2849400, 2851200, 2853000, 2854800, 
    2856600, 2858400, 2860200, 2862000, 2863800, 2865600, 2867400, 2869200, 
    2871000, 2872800, 2874600, 2876400, 2878200, 2880000, 2881800, 2883600, 
    2885400, 2887200, 2889000, 2890800, 2892600, 2894400, 2896200, 2898000, 
    2899800, 2901600, 2903400, 2905200, 2907000, 2908800, 2910600, 2912400, 
    2914200, 2916000, 2917800, 2919600, 2921400, 2923200, 2925000, 2926800, 
    2928600, 2930400, 2932200, 2934000, 2935800, 2937600, 2939400, 2941200, 
    2943000, 2944800, 2946600, 2948400, 2950200, 2952000, 2953800, 2955600, 
    2957400, 2959200, 2961000, 2962800, 2964600, 2966400, 2968200, 2970000, 
    2971800, 2973600, 2975400, 2977200, 2979000, 2980800, 2982600, 2984400, 
    2986200, 2988000, 2989800, 2991600, 2993400, 2995200, 2997000, 2998800, 
    3000600, 3002400, 3004200, 3006000, 3007800, 3009600, 3011400, 3013200, 
    3015000, 3016800, 3018600, 3020400, 3022200, 3024000, 3025800, 3027600, 
    3029400, 3031200, 3033000, 3034800, 3036600, 3038400, 3040200, 3042000, 
    3043800, 3045600, 3047400, 3049200, 3051000, 3052800, 3054600, 3056400, 
    3058200, 3060000, 3061800, 3063600, 3065400, 3067200, 3069000, 3070800, 
    3072600, 3074400, 3076200, 3078000, 3079800, 3081600, 3083400, 3085200, 
    3087000, 3088800, 3090600, 3092400, 3094200, 3096000, 3097800, 3099600, 
    3101400, 3103200, 3105000, 3106800, 3108600, 3110400, 3112200, 3114000, 
    3115800, 3117600, 3119400, 3121200, 3123000, 3124800, 3126600, 3128400, 
    3130200, 3132000, 3133800, 3135600, 3137400, 3139200, 3141000, 3142800, 
    3144600, 3146400, 3148200, 3150000, 3151800, 3153600, 3155400, 3157200, 
    3159000, 3160800, 3162600, 3164400, 3166200, 3168000, 3169800, 3171600, 
    3173400, 3175200, 3177000, 3178800, 3180600, 3182400, 3184200, 3186000, 
    3187800, 3189600, 3191400, 3193200, 3195000, 3196800, 3198600, 3200400, 
    3202200, 3204000, 3205800, 3207600, 3209400, 3211200, 3213000, 3214800, 
    3216600, 3218400, 3220200, 3222000, 3223800, 3225600, 3227400, 3229200, 
    3231000, 3232800, 3234600, 3236400, 3238200, 3240000, 3241800, 3243600, 
    3245400, 3247200, 3249000, 3250800, 3252600, 3254400, 3256200, 3258000, 
    3259800, 3261600, 3263400, 3265200, 3267000, 3268800, 3270600, 3272400, 
    3274200, 3276000, 3277800, 3279600, 3281400, 3283200, 3285000, 3286800, 
    3288600, 3290400, 3292200, 3294000, 3295800, 3297600, 3299400, 3301200, 
    3303000, 3304800, 3306600, 3308400, 3310200, 3312000, 3313800, 3315600, 
    3317400, 3319200, 3321000, 3322800, 3324600, 3326400, 3328200, 3330000, 
    3331800, 3333600, 3335400, 3337200, 3339000, 3340800, 3342600, 3344400, 
    3346200, 3348000, 3349800, 3351600, 3353400, 3355200, 3357000, 3358800, 
    3360600, 3362400, 3364200, 3366000, 3367800, 3369600, 3371400, 3373200, 
    3375000, 3376800, 3378600, 3380400, 3382200, 3384000, 3385800, 3387600, 
    3389400, 3391200, 3393000, 3394800, 3396600, 3398400, 3400200, 3402000, 
    3403800, 3405600, 3407400, 3409200, 3411000, 3412800, 3414600, 3416400, 
    3418200, 3420000, 3421800, 3423600, 3425400, 3427200, 3429000, 3430800, 
    3432600, 3434400, 3436200, 3438000, 3439800, 3441600, 3443400, 3445200, 
    3447000, 3448800, 3450600, 3452400, 3454200, 3456000, 3457800, 3459600, 
    3461400, 3463200, 3465000, 3466800, 3468600, 3470400, 3472200, 3474000, 
    3475800, 3477600, 3479400, 3481200, 3483000, 3484800, 3486600, 3488400, 
    3490200, 3492000, 3493800, 3495600, 3497400, 3499200, 3501000, 3502800, 
    3504600, 3506400, 3508200, 3510000, 3511800, 3513600, 3515400, 3517200, 
    3519000, 3520800, 3522600, 3524400, 3526200, 3528000, 3529800, 3531600, 
    3533400, 3535200, 3537000, 3538800, 3540600, 3542400, 3544200, 3546000, 
    3547800, 3549600, 3551400, 3553200, 3555000, 3556800, 3558600, 3560400, 
    3562200, 3564000, 3565800, 3567600, 3569400, 3571200, 3573000, 3574800, 
    3576600, 3578400, 3580200, 3582000, 3583800, 3585600, 3587400, 3589200, 
    3591000, 3592800, 3594600, 3596400, 3598200, 3600000, 3601800, 3603600, 
    3605400, 3607200, 3609000, 3610800, 3612600, 3614400, 3616200, 3618000, 
    3619800, 3621600, 3623400, 3625200, 3627000, 3628800, 3630600, 3632400, 
    3634200, 3636000, 3637800, 3639600, 3641400, 3643200, 3645000, 3646800, 
    3648600, 3650400, 3652200, 3654000, 3655800, 3657600, 3659400, 3661200, 
    3663000, 3664800, 3666600, 3668400, 3670200, 3672000, 3673800, 3675600, 
    3677400, 3679200, 3681000, 3682800, 3684600, 3686400, 3688200, 3690000, 
    3691800, 3693600, 3695400, 3697200, 3699000, 3700800, 3702600, 3704400, 
    3706200, 3708000, 3709800, 3711600, 3713400, 3715200, 3717000, 3718800, 
    3720600, 3722400, 3724200, 3726000, 3727800, 3729600, 3731400, 3733200, 
    3735000, 3736800, 3738600, 3740400, 3742200, 3744000, 3745800, 3747600, 
    3749400, 3751200, 3753000, 3754800, 3756600, 3758400, 3760200, 3762000, 
    3763800, 3765600, 3767400, 3769200, 3771000, 3772800, 3774600, 3776400, 
    3778200, 3780000, 3781800, 3783600, 3785400, 3787200, 3789000, 3790800, 
    3792600, 3794400, 3796200, 3798000, 3799800, 3801600, 3803400, 3805200, 
    3807000, 3808800, 3810600, 3812400, 3814200, 3816000, 3817800, 3819600, 
    3821400, 3823200, 3825000, 3826800, 3828600, 3830400, 3832200, 3834000, 
    3835800, 3837600, 3839400, 3841200, 3843000, 3844800, 3846600, 3848400, 
    3850200, 3852000, 3853800, 3855600, 3857400, 3859200, 3861000, 3862800, 
    3864600, 3866400, 3868200, 3870000, 3871800, 3873600, 3875400, 3877200, 
    3879000, 3880800, 3882600, 3884400, 3886200, 3888000, 3889800, 3891600, 
    3893400, 3895200, 3897000, 3898800, 3900600, 3902400, 3904200, 3906000, 
    3907800, 3909600, 3911400, 3913200, 3915000, 3916800, 3918600, 3920400, 
    3922200, 3924000, 3925800, 3927600, 3929400, 3931200, 3933000, 3934800, 
    3936600, 3938400, 3940200, 3942000, 3943800, 3945600, 3947400, 3949200, 
    3951000, 3952800, 3954600, 3956400, 3958200, 3960000, 3961800, 3963600, 
    3965400, 3967200, 3969000, 3970800, 3972600, 3974400, 3976200, 3978000, 
    3979800, 3981600, 3983400, 3985200, 3987000, 3988800, 3990600, 3992400, 
    3994200, 3996000, 3997800, 3999600, 4001400, 4003200, 4005000, 4006800, 
    4008600, 4010400, 4012200, 4014000, 4015800, 4017600, 4019400, 4021200, 
    4023000, 4024800, 4026600, 4028400, 4030200, 4032000, 4033800, 4035600, 
    4037400, 4039200, 4041000, 4042800, 4044600, 4046400, 4048200, 4050000, 
    4051800, 4053600, 4055400, 4057200, 4059000, 4060800, 4062600, 4064400, 
    4066200, 4068000, 4069800, 4071600, 4073400, 4075200, 4077000, 4078800, 
    4080600, 4082400, 4084200, 4086000, 4087800, 4089600, 4091400, 4093200, 
    4095000, 4096800, 4098600, 4100400, 4102200, 4104000, 4105800, 4107600, 
    4109400, 4111200, 4113000, 4114800, 4116600, 4118400, 4120200, 4122000, 
    4123800, 4125600, 4127400, 4129200, 4131000, 4132800, 4134600, 4136400, 
    4138200, 4140000, 4141800, 4143600, 4145400, 4147200, 4149000, 4150800, 
    4152600, 4154400, 4156200, 4158000, 4159800, 4161600, 4163400, 4165200, 
    4167000, 4168800, 4170600, 4172400, 4174200, 4176000, 4177800, 4179600, 
    4181400, 4183200, 4185000, 4186800, 4188600, 4190400, 4192200, 4194000, 
    4195800, 4197600, 4199400, 4201200, 4203000, 4204800, 4206600, 4208400, 
    4210200, 4212000, 4213800, 4215600, 4217400, 4219200, 4221000, 4222800, 
    4224600, 4226400, 4228200, 4230000, 4231800, 4233600, 4235400, 4237200, 
    4239000, 4240800, 4242600, 4244400, 4246200, 4248000, 4249800, 4251600, 
    4253400, 4255200, 4257000, 4258800, 4260600, 4262400, 4264200, 4266000, 
    4267800, 4269600, 4271400, 4273200, 4275000, 4276800, 4278600, 4280400, 
    4282200, 4284000, 4285800, 4287600, 4289400, 4291200, 4293000, 4294800, 
    4296600, 4298400, 4300200, 4302000, 4303800, 4305600, 4307400, 4309200, 
    4311000, 4312800, 4314600, 4316400, 4318200, 4320000, 4321800, 4323600, 
    4325400, 4327200, 4329000, 4330800, 4332600, 4334400, 4336200, 4338000, 
    4339800, 4341600, 4343400, 4345200, 4347000, 4348800, 4350600, 4352400, 
    4354200, 4356000, 4357800, 4359600, 4361400, 4363200, 4365000, 4366800, 
    4368600, 4370400, 4372200, 4374000, 4375800, 4377600, 4379400, 4381200, 
    4383000, 4384800, 4386600, 4388400, 4390200, 4392000, 4393800, 4395600, 
    4397400, 4399200, 4401000, 4402800, 4404600, 4406400, 4408200, 4410000, 
    4411800, 4413600, 4415400, 4417200, 4419000, 4420800, 4422600, 4424400, 
    4426200, 4428000, 4429800, 4431600, 4433400, 4435200, 4437000, 4438800, 
    4440600, 4442400, 4444200, 4446000, 4447800, 4449600, 4451400, 4453200, 
    4455000, 4456800, 4458600, 4460400, 4462200, 4464000, 4465800, 4467600, 
    4469400, 4471200, 4473000, 4474800, 4476600, 4478400, 4480200, 4482000, 
    4483800, 4485600, 4487400, 4489200, 4491000, 4492800, 4494600, 4496400, 
    4498200, 4500000, 4501800, 4503600, 4505400, 4507200, 4509000, 4510800, 
    4512600, 4514400, 4516200, 4518000, 4519800, 4521600, 4523400, 4525200, 
    4527000, 4528800, 4530600, 4532400, 4534200, 4536000, 4537800, 4539600, 
    4541400, 4543200, 4545000, 4546800, 4548600, 4550400, 4552200, 4554000, 
    4555800, 4557600, 4559400, 4561200, 4563000, 4564800, 4566600, 4568400, 
    4570200, 4572000, 4573800, 4575600, 4577400, 4579200, 4581000, 4582800, 
    4584600, 4586400, 4588200, 4590000, 4591800, 4593600, 4595400, 4597200, 
    4599000, 4600800, 4602600, 4604400, 4606200, 4608000, 4609800, 4611600, 
    4613400, 4615200, 4617000, 4618800, 4620600, 4622400, 4624200, 4626000, 
    4627800, 4629600, 4631400, 4633200, 4635000, 4636800, 4638600, 4640400, 
    4642200, 4644000, 4645800, 4647600, 4649400, 4651200, 4653000, 4654800, 
    4656600, 4658400, 4660200, 4662000, 4663800, 4665600, 4667400, 4669200, 
    4671000, 4672800, 4674600, 4676400, 4678200, 4680000, 4681800, 4683600, 
    4685400, 4687200, 4689000, 4690800, 4692600, 4694400, 4696200, 4698000, 
    4699800, 4701600, 4703400, 4705200, 4707000, 4708800, 4710600, 4712400, 
    4714200, 4716000, 4717800, 4719600, 4721400, 4723200, 4725000, 4726800, 
    4728600, 4730400, 4732200, 4734000, 4735800, 4737600, 4739400, 4741200, 
    4743000, 4744800, 4746600, 4748400, 4750200, 4752000, 4753800, 4755600, 
    4757400, 4759200, 4761000, 4762800, 4764600, 4766400, 4768200, 4770000, 
    4771800, 4773600, 4775400, 4777200, 4779000, 4780800, 4782600, 4784400, 
    4786200, 4788000, 4789800, 4791600, 4793400, 4795200, 4797000, 4798800, 
    4800600, 4802400, 4804200, 4806000, 4807800, 4809600, 4811400, 4813200, 
    4815000, 4816800, 4818600, 4820400, 4822200, 4824000, 4825800, 4827600, 
    4829400, 4831200, 4833000, 4834800, 4836600, 4838400, 4840200, 4842000, 
    4843800, 4845600, 4847400, 4849200, 4851000, 4852800, 4854600, 4856400, 
    4858200, 4860000, 4861800, 4863600, 4865400, 4867200, 4869000, 4870800, 
    4872600, 4874400, 4876200, 4878000, 4879800, 4881600, 4883400, 4885200, 
    4887000, 4888800, 4890600, 4892400, 4894200, 4896000, 4897800, 4899600, 
    4901400, 4903200, 4905000, 4906800, 4908600, 4910400, 4912200, 4914000, 
    4915800, 4917600, 4919400, 4921200, 4923000, 4924800, 4926600, 4928400, 
    4930200, 4932000, 4933800, 4935600, 4937400, 4939200, 4941000, 4942800, 
    4944600, 4946400, 4948200, 4950000, 4951800, 4953600, 4955400, 4957200, 
    4959000, 4960800, 4962600, 4964400, 4966200, 4968000, 4969800, 4971600, 
    4973400, 4975200, 4977000, 4978800, 4980600, 4982400, 4984200, 4986000, 
    4987800, 4989600, 4991400, 4993200, 4995000, 4996800, 4998600, 5000400, 
    5002200, 5004000, 5005800, 5007600, 5009400, 5011200, 5013000, 5014800, 
    5016600, 5018400, 5020200, 5022000, 5023800, 5025600, 5027400, 5029200, 
    5031000, 5032800, 5034600, 5036400, 5038200, 5040000, 5041800, 5043600, 
    5045400, 5047200, 5049000, 5050800, 5052600, 5054400, 5056200, 5058000, 
    5059800, 5061600, 5063400, 5065200, 5067000, 5068800, 5070600, 5072400, 
    5074200, 5076000, 5077800, 5079600, 5081400, 5083200, 5085000, 5086800, 
    5088600, 5090400, 5092200, 5094000, 5095800, 5097600, 5099400, 5101200, 
    5103000, 5104800, 5106600, 5108400, 5110200, 5112000, 5113800, 5115600, 
    5117400, 5119200, 5121000, 5122800, 5124600, 5126400, 5128200, 5130000, 
    5131800, 5133600, 5135400, 5137200, 5139000, 5140800, 5142600, 5144400, 
    5146200, 5148000, 5149800, 5151600, 5153400, 5155200, 5157000, 5158800, 
    5160600, 5162400, 5164200, 5166000, 5167800, 5169600, 5171400, 5173200, 
    5175000, 5176800, 5178600, 5180400, 5182200, 5184000, 5185800, 5187600, 
    5189400, 5191200, 5193000, 5194800, 5196600, 5198400, 5200200, 5202000, 
    5203800, 5205600, 5207400, 5209200, 5211000, 5212800, 5214600, 5216400, 
    5218200, 5220000, 5221800, 5223600, 5225400, 5227200, 5229000, 5230800, 
    5232600, 5234400, 5236200, 5238000, 5239800, 5241600, 5243400, 5245200, 
    5247000, 5248800, 5250600, 5252400, 5254200, 5256000, 5257800, 5259600, 
    5261400, 5263200, 5265000, 5266800, 5268600, 5270400, 5272200, 5274000, 
    5275800, 5277600, 5279400, 5281200, 5283000, 5284800, 5286600, 5288400, 
    5290200, 5292000, 5293800, 5295600, 5297400, 5299200, 5301000, 5302800, 
    5304600, 5306400, 5308200, 5310000, 5311800, 5313600, 5315400, 5317200, 
    5319000, 5320800, 5322600, 5324400, 5326200, 5328000, 5329800, 5331600, 
    5333400, 5335200, 5337000, 5338800, 5340600, 5342400, 5344200, 5346000, 
    5347800, 5349600, 5351400, 5353200, 5355000, 5356800, 5358600, 5360400, 
    5362200, 5364000, 5365800, 5367600, 5369400, 5371200, 5373000, 5374800, 
    5376600, 5378400, 5380200, 5382000, 5383800, 5385600, 5387400, 5389200, 
    5391000, 5392800, 5394600, 5396400, 5398200, 5400000, 5401800, 5403600, 
    5405400, 5407200, 5409000, 5410800, 5412600, 5414400, 5416200, 5418000, 
    5419800, 5421600, 5423400, 5425200, 5427000, 5428800, 5430600, 5432400, 
    5434200, 5436000, 5437800, 5439600, 5441400, 5443200, 5445000, 5446800, 
    5448600, 5450400, 5452200, 5454000, 5455800, 5457600, 5459400, 5461200, 
    5463000, 5464800, 5466600, 5468400, 5470200, 5472000, 5473800, 5475600, 
    5477400, 5479200, 5481000, 5482800, 5484600, 5486400, 5488200, 5490000, 
    5491800, 5493600, 5495400, 5497200, 5499000, 5500800, 5502600, 5504400, 
    5506200, 5508000, 5509800, 5511600, 5513400, 5515200, 5517000, 5518800, 
    5520600, 5522400, 5524200, 5526000, 5527800, 5529600, 5531400, 5533200, 
    5535000, 5536800, 5538600, 5540400, 5542200, 5544000, 5545800, 5547600, 
    5549400, 5551200, 5553000, 5554800, 5556600, 5558400, 5560200, 5562000, 
    5563800, 5565600, 5567400, 5569200, 5571000, 5572800, 5574600, 5576400, 
    5578200, 5580000, 5581800, 5583600, 5585400, 5587200, 5589000, 5590800, 
    5592600, 5594400, 5596200, 5598000, 5599800, 5601600, 5603400, 5605200, 
    5607000, 5608800, 5610600, 5612400, 5614200, 5616000, 5617800, 5619600, 
    5621400, 5623200, 5625000, 5626800, 5628600, 5630400, 5632200, 5634000, 
    5635800, 5637600, 5639400, 5641200, 5643000, 5644800, 5646600, 5648400, 
    5650200, 5652000, 5653800, 5655600, 5657400, 5659200, 5661000, 5662800, 
    5664600, 5666400, 5668200, 5670000, 5671800, 5673600, 5675400, 5677200, 
    5679000, 5680800, 5682600, 5684400, 5686200, 5688000, 5689800, 5691600, 
    5693400, 5695200, 5697000, 5698800, 5700600, 5702400, 5704200, 5706000, 
    5707800, 5709600, 5711400, 5713200, 5715000, 5716800, 5718600, 5720400, 
    5722200, 5724000, 5725800, 5727600, 5729400, 5731200, 5733000, 5734800, 
    5736600, 5738400, 5740200, 5742000, 5743800, 5745600, 5747400, 5749200, 
    5751000, 5752800, 5754600, 5756400, 5758200, 5760000, 5761800, 5763600, 
    5765400, 5767200, 5769000, 5770800, 5772600, 5774400, 5776200, 5778000, 
    5779800, 5781600, 5783400, 5785200, 5787000, 5788800, 5790600, 5792400, 
    5794200, 5796000, 5797800, 5799600, 5801400, 5803200, 5805000, 5806800, 
    5808600, 5810400, 5812200, 5814000, 5815800, 5817600, 5819400, 5821200, 
    5823000, 5824800, 5826600, 5828400, 5830200, 5832000, 5833800, 5835600, 
    5837400, 5839200, 5841000, 5842800, 5844600, 5846400, 5848200, 5850000, 
    5851800, 5853600, 5855400, 5857200, 5859000, 5860800, 5862600, 5864400, 
    5866200, 5868000, 5869800, 5871600, 5873400, 5875200, 5877000, 5878800, 
    5880600, 5882400, 5884200, 5886000, 5887800, 5889600, 5891400, 5893200, 
    5895000, 5896800, 5898600, 5900400, 5902200, 5904000, 5905800, 5907600, 
    5909400, 5911200, 5913000, 5914800, 5916600, 5918400, 5920200, 5922000, 
    5923800, 5925600, 5927400, 5929200, 5931000, 5932800, 5934600, 5936400, 
    5938200, 5940000, 5941800, 5943600, 5945400, 5947200, 5949000, 5950800, 
    5952600, 5954400, 5956200, 5958000, 5959800, 5961600, 5963400, 5965200, 
    5967000, 5968800, 5970600, 5972400, 5974200, 5976000, 5977800, 5979600, 
    5981400, 5983200, 5985000, 5986800, 5988600, 5990400, 5992200, 5994000, 
    5995800, 5997600, 5999400, 6001200, 6003000, 6004800, 6006600, 6008400, 
    6010200, 6012000, 6013800, 6015600, 6017400, 6019200, 6021000, 6022800, 
    6024600, 6026400, 6028200, 6030000, 6031800, 6033600, 6035400, 6037200, 
    6039000, 6040800, 6042600, 6044400, 6046200, 6048000, 6049800, 6051600, 
    6053400, 6055200, 6057000, 6058800, 6060600, 6062400, 6064200, 6066000, 
    6067800, 6069600, 6071400, 6073200, 6075000, 6076800, 6078600, 6080400, 
    6082200, 6084000, 6085800, 6087600, 6089400, 6091200, 6093000, 6094800, 
    6096600, 6098400, 6100200, 6102000, 6103800, 6105600, 6107400, 6109200, 
    6111000, 6112800, 6114600, 6116400, 6118200, 6120000, 6121800, 6123600, 
    6125400, 6127200, 6129000, 6130800, 6132600, 6134400, 6136200, 6138000, 
    6139800, 6141600, 6143400, 6145200, 6147000, 6148800, 6150600, 6152400, 
    6154200, 6156000, 6157800, 6159600, 6161400, 6163200, 6165000, 6166800, 
    6168600, 6170400, 6172200, 6174000, 6175800, 6177600, 6179400, 6181200, 
    6183000, 6184800, 6186600, 6188400, 6190200, 6192000, 6193800, 6195600, 
    6197400, 6199200, 6201000, 6202800, 6204600, 6206400, 6208200, 6210000, 
    6211800, 6213600, 6215400, 6217200, 6219000, 6220800, 6222600, 6224400, 
    6226200, 6228000, 6229800, 6231600, 6233400, 6235200, 6237000, 6238800, 
    6240600, 6242400, 6244200, 6246000, 6247800, 6249600, 6251400, 6253200, 
    6255000, 6256800, 6258600, 6260400, 6262200, 6264000, 6265800, 6267600, 
    6269400, 6271200, 6273000, 6274800, 6276600, 6278400, 6280200, 6282000, 
    6283800, 6285600, 6287400, 6289200, 6291000, 6292800, 6294600, 6296400, 
    6298200, 6300000, 6301800, 6303600, 6305400, 6307200, 6309000, 6310800, 
    6312600, 6314400, 6316200, 6318000, 6319800, 6321600, 6323400, 6325200, 
    6327000, 6328800, 6330600, 6332400, 6334200, 6336000, 6337800, 6339600, 
    6341400, 6343200, 6345000, 6346800, 6348600, 6350400, 6352200, 6354000, 
    6355800, 6357600, 6359400, 6361200, 6363000, 6364800, 6366600, 6368400, 
    6370200, 6372000, 6373800, 6375600, 6377400, 6379200, 6381000, 6382800, 
    6384600, 6386400, 6388200, 6390000, 6391800, 6393600, 6395400, 6397200, 
    6399000, 6400800, 6402600, 6404400, 6406200, 6408000, 6409800, 6411600, 
    6413400, 6415200, 6417000, 6418800, 6420600, 6422400, 6424200, 6426000, 
    6427800, 6429600, 6431400, 6433200, 6435000, 6436800, 6438600, 6440400, 
    6442200, 6444000, 6445800, 6447600, 6449400, 6451200, 6453000, 6454800, 
    6456600, 6458400, 6460200, 6462000, 6463800, 6465600, 6467400, 6469200, 
    6471000, 6472800, 6474600, 6476400, 6478200, 6480000, 6481800, 6483600, 
    6485400, 6487200, 6489000, 6490800, 6492600, 6494400, 6496200, 6498000, 
    6499800, 6501600, 6503400, 6505200, 6507000, 6508800, 6510600, 6512400, 
    6514200, 6516000, 6517800, 6519600, 6521400, 6523200, 6525000, 6526800, 
    6528600, 6530400, 6532200, 6534000, 6535800, 6537600, 6539400, 6541200, 
    6543000, 6544800, 6546600, 6548400, 6550200, 6552000, 6553800, 6555600, 
    6557400, 6559200, 6561000, 6562800, 6564600, 6566400, 6568200, 6570000, 
    6571800, 6573600, 6575400, 6577200, 6579000, 6580800, 6582600, 6584400, 
    6586200, 6588000, 6589800, 6591600, 6593400, 6595200, 6597000, 6598800, 
    6600600, 6602400, 6604200, 6606000, 6607800, 6609600, 6611400, 6613200, 
    6615000, 6616800, 6618600, 6620400, 6622200, 6624000, 6625800, 6627600, 
    6629400, 6631200, 6633000, 6634800, 6636600, 6638400, 6640200, 6642000, 
    6643800, 6645600, 6647400, 6649200, 6651000, 6652800, 6654600, 6656400, 
    6658200, 6660000, 6661800, 6663600, 6665400, 6667200, 6669000, 6670800, 
    6672600, 6674400, 6676200, 6678000, 6679800, 6681600, 6683400, 6685200, 
    6687000, 6688800, 6690600, 6692400, 6694200, 6696000, 6697800, 6699600, 
    6701400, 6703200, 6705000, 6706800, 6708600, 6710400, 6712200, 6714000, 
    6715800, 6717600, 6719400, 6721200, 6723000, 6724800, 6726600, 6728400, 
    6730200, 6732000, 6733800, 6735600, 6737400, 6739200, 6741000, 6742800, 
    6744600, 6746400, 6748200, 6750000, 6751800, 6753600, 6755400, 6757200, 
    6759000, 6760800, 6762600, 6764400, 6766200, 6768000, 6769800, 6771600, 
    6773400, 6775200, 6777000, 6778800, 6780600, 6782400, 6784200, 6786000, 
    6787800, 6789600, 6791400, 6793200, 6795000, 6796800, 6798600, 6800400, 
    6802200, 6804000, 6805800, 6807600, 6809400, 6811200, 6813000, 6814800, 
    6816600, 6818400, 6820200, 6822000, 6823800, 6825600, 6827400, 6829200, 
    6831000, 6832800, 6834600, 6836400, 6838200, 6840000, 6841800, 6843600, 
    6845400, 6847200, 6849000, 6850800, 6852600, 6854400, 6856200, 6858000, 
    6859800, 6861600, 6863400, 6865200, 6867000, 6868800, 6870600, 6872400, 
    6874200, 6876000, 6877800, 6879600, 6881400, 6883200, 6885000, 6886800, 
    6888600, 6890400, 6892200, 6894000, 6895800, 6897600, 6899400, 6901200, 
    6903000, 6904800, 6906600, 6908400, 6910200, 6912000, 6913800, 6915600, 
    6917400, 6919200, 6921000, 6922800, 6924600, 6926400, 6928200, 6930000, 
    6931800, 6933600, 6935400, 6937200, 6939000, 6940800, 6942600, 6944400, 
    6946200, 6948000, 6949800, 6951600, 6953400, 6955200, 6957000, 6958800, 
    6960600, 6962400, 6964200, 6966000, 6967800, 6969600, 6971400, 6973200, 
    6975000, 6976800, 6978600, 6980400, 6982200, 6984000, 6985800, 6987600, 
    6989400, 6991200, 6993000, 6994800, 6996600, 6998400, 7000200, 7002000, 
    7003800, 7005600, 7007400, 7009200, 7011000, 7012800, 7014600, 7016400, 
    7018200, 7020000, 7021800, 7023600, 7025400, 7027200, 7029000, 7030800, 
    7032600, 7034400, 7036200, 7038000, 7039800, 7041600, 7043400, 7045200, 
    7047000, 7048800, 7050600, 7052400, 7054200, 7056000, 7057800, 7059600, 
    7061400, 7063200, 7065000, 7066800, 7068600, 7070400, 7072200, 7074000, 
    7075800, 7077600, 7079400, 7081200, 7083000, 7084800, 7086600, 7088400, 
    7090200, 7092000, 7093800, 7095600, 7097400, 7099200, 7101000, 7102800, 
    7104600, 7106400, 7108200, 7110000, 7111800, 7113600, 7115400, 7117200, 
    7119000, 7120800, 7122600, 7124400, 7126200, 7128000, 7129800, 7131600, 
    7133400, 7135200, 7137000, 7138800, 7140600, 7142400, 7144200, 7146000, 
    7147800, 7149600, 7151400, 7153200, 7155000, 7156800, 7158600, 7160400, 
    7162200, 7164000, 7165800, 7167600, 7169400, 7171200, 7173000, 7174800, 
    7176600, 7178400, 7180200, 7182000, 7183800, 7185600, 7187400, 7189200, 
    7191000, 7192800, 7194600, 7196400, 7198200, 7200000, 7201800, 7203600, 
    7205400, 7207200, 7209000, 7210800, 7212600, 7214400, 7216200, 7218000, 
    7219800, 7221600, 7223400, 7225200, 7227000, 7228800, 7230600, 7232400, 
    7234200, 7236000, 7237800, 7239600, 7241400, 7243200, 7245000, 7246800, 
    7248600, 7250400, 7252200, 7254000, 7255800, 7257600, 7259400, 7261200, 
    7263000, 7264800, 7266600, 7268400, 7270200, 7272000, 7273800, 7275600, 
    7277400, 7279200, 7281000, 7282800, 7284600, 7286400, 7288200, 7290000, 
    7291800, 7293600, 7295400, 7297200, 7299000, 7300800, 7302600, 7304400, 
    7306200, 7308000, 7309800, 7311600, 7313400, 7315200, 7317000, 7318800, 
    7320600, 7322400, 7324200, 7326000, 7327800, 7329600, 7331400, 7333200, 
    7335000, 7336800, 7338600, 7340400, 7342200, 7344000, 7345800, 7347600, 
    7349400, 7351200, 7353000, 7354800, 7356600, 7358400, 7360200, 7362000, 
    7363800, 7365600, 7367400, 7369200, 7371000, 7372800, 7374600, 7376400, 
    7378200, 7380000, 7381800, 7383600, 7385400, 7387200, 7389000, 7390800, 
    7392600, 7394400, 7396200, 7398000, 7399800, 7401600, 7403400, 7405200, 
    7407000, 7408800, 7410600, 7412400, 7414200, 7416000, 7417800, 7419600, 
    7421400, 7423200, 7425000, 7426800, 7428600, 7430400, 7432200, 7434000, 
    7435800, 7437600, 7439400, 7441200, 7443000, 7444800, 7446600, 7448400, 
    7450200, 7452000, 7453800, 7455600, 7457400, 7459200, 7461000, 7462800, 
    7464600, 7466400, 7468200, 7470000, 7471800, 7473600, 7475400, 7477200, 
    7479000, 7480800, 7482600, 7484400, 7486200, 7488000, 7489800, 7491600, 
    7493400, 7495200, 7497000, 7498800, 7500600, 7502400, 7504200, 7506000, 
    7507800, 7509600, 7511400, 7513200, 7515000, 7516800, 7518600, 7520400, 
    7522200, 7524000, 7525800, 7527600, 7529400, 7531200, 7533000, 7534800, 
    7536600, 7538400, 7540200, 7542000, 7543800, 7545600, 7547400, 7549200, 
    7551000, 7552800, 7554600, 7556400, 7558200, 7560000, 7561800, 7563600, 
    7565400, 7567200, 7569000, 7570800, 7572600, 7574400, 7576200, 7578000, 
    7579800, 7581600, 7583400, 7585200, 7587000, 7588800, 7590600, 7592400, 
    7594200, 7596000, 7597800, 7599600, 7601400, 7603200, 7605000, 7606800, 
    7608600, 7610400, 7612200, 7614000, 7615800, 7617600, 7619400, 7621200, 
    7623000, 7624800, 7626600, 7628400, 7630200, 7632000, 7633800, 7635600, 
    7637400, 7639200, 7641000, 7642800, 7644600, 7646400, 7648200, 7650000, 
    7651800, 7653600, 7655400, 7657200, 7659000, 7660800, 7662600, 7664400, 
    7666200, 7668000, 7669800, 7671600, 7673400, 7675200, 7677000, 7678800, 
    7680600, 7682400, 7684200, 7686000, 7687800, 7689600, 7691400, 7693200, 
    7695000, 7696800, 7698600, 7700400, 7702200, 7704000, 7705800, 7707600, 
    7709400, 7711200, 7713000, 7714800, 7716600, 7718400, 7720200, 7722000, 
    7723800, 7725600, 7727400, 7729200, 7731000, 7732800, 7734600, 7736400, 
    7738200, 7740000, 7741800, 7743600, 7745400, 7747200, 7749000, 7750800, 
    7752600, 7754400, 7756200, 7758000, 7759800, 7761600, 7763400, 7765200, 
    7767000, 7768800, 7770600, 7772400, 7774200, 7776000, 7777800, 7779600, 
    7781400, 7783200, 7785000, 7786800, 7788600, 7790400, 7792200, 7794000, 
    7795800, 7797600, 7799400, 7801200, 7803000, 7804800, 7806600, 7808400, 
    7810200, 7812000, 7813800, 7815600, 7817400, 7819200, 7821000, 7822800, 
    7824600, 7826400, 7828200, 7830000, 7831800, 7833600, 7835400, 7837200, 
    7839000, 7840800, 7842600, 7844400, 7846200, 7848000, 7849800, 7851600, 
    7853400, 7855200, 7857000, 7858800, 7860600, 7862400, 7864200, 7866000, 
    7867800, 7869600, 7871400, 7873200, 7875000, 7876800, 7878600, 7880400, 
    7882200, 7884000, 7885800, 7887600, 7889400, 7891200, 7893000, 7894800, 
    7896600, 7898400, 7900200, 7902000, 7903800, 7905600, 7907400, 7909200, 
    7911000, 7912800, 7914600, 7916400, 7918200, 7920000, 7921800, 7923600, 
    7925400, 7927200, 7929000, 7930800, 7932600, 7934400, 7936200, 7938000, 
    7939800, 7941600, 7943400, 7945200, 7947000, 7948800, 7950600, 7952400, 
    7954200, 7956000, 7957800, 7959600, 7961400, 7963200, 7965000, 7966800, 
    7968600, 7970400, 7972200, 7974000, 7975800, 7977600, 7979400, 7981200, 
    7983000, 7984800, 7986600, 7988400, 7990200, 7992000, 7993800, 7995600, 
    7997400, 7999200, 8001000, 8002800, 8004600, 8006400, 8008200, 8010000, 
    8011800, 8013600, 8015400, 8017200, 8019000, 8020800, 8022600, 8024400, 
    8026200, 8028000, 8029800, 8031600, 8033400, 8035200, 8037000, 8038800, 
    8040600, 8042400, 8044200, 8046000, 8047800, 8049600, 8051400, 8053200, 
    8055000, 8056800, 8058600, 8060400, 8062200, 8064000, 8065800, 8067600, 
    8069400, 8071200, 8073000, 8074800, 8076600, 8078400, 8080200, 8082000, 
    8083800, 8085600, 8087400, 8089200, 8091000, 8092800, 8094600, 8096400, 
    8098200, 8100000, 8101800, 8103600, 8105400, 8107200, 8109000, 8110800, 
    8112600, 8114400, 8116200, 8118000, 8119800, 8121600, 8123400, 8125200, 
    8127000, 8128800, 8130600, 8132400, 8134200, 8136000, 8137800, 8139600, 
    8141400, 8143200, 8145000, 8146800, 8148600, 8150400, 8152200, 8154000, 
    8155800, 8157600, 8159400, 8161200, 8163000, 8164800, 8166600, 8168400, 
    8170200, 8172000, 8173800, 8175600, 8177400, 8179200, 8181000, 8182800, 
    8184600, 8186400, 8188200, 8190000, 8191800, 8193600, 8195400, 8197200, 
    8199000, 8200800, 8202600, 8204400, 8206200, 8208000, 8209800, 8211600, 
    8213400, 8215200, 8217000, 8218800, 8220600, 8222400, 8224200, 8226000, 
    8227800, 8229600, 8231400, 8233200, 8235000, 8236800, 8238600, 8240400, 
    8242200, 8244000, 8245800, 8247600, 8249400, 8251200, 8253000, 8254800, 
    8256600, 8258400, 8260200, 8262000, 8263800, 8265600, 8267400, 8269200, 
    8271000, 8272800, 8274600, 8276400, 8278200, 8280000, 8281800, 8283600, 
    8285400, 8287200, 8289000, 8290800, 8292600, 8294400, 8296200, 8298000, 
    8299800, 8301600, 8303400, 8305200, 8307000, 8308800, 8310600, 8312400, 
    8314200, 8316000, 8317800, 8319600, 8321400, 8323200, 8325000, 8326800, 
    8328600, 8330400, 8332200, 8334000, 8335800, 8337600, 8339400, 8341200, 
    8343000, 8344800, 8346600, 8348400, 8350200, 8352000, 8353800, 8355600, 
    8357400, 8359200, 8361000, 8362800, 8364600, 8366400, 8368200, 8370000, 
    8371800, 8373600, 8375400, 8377200, 8379000, 8380800, 8382600, 8384400, 
    8386200, 8388000, 8389800, 8391600, 8393400, 8395200, 8397000, 8398800, 
    8400600, 8402400, 8404200, 8406000, 8407800, 8409600, 8411400, 8413200, 
    8415000, 8416800, 8418600, 8420400, 8422200, 8424000, 8425800, 8427600, 
    8429400, 8431200, 8433000, 8434800, 8436600, 8438400, 8440200, 8442000, 
    8443800, 8445600, 8447400, 8449200, 8451000, 8452800, 8454600, 8456400, 
    8458200, 8460000, 8461800, 8463600, 8465400, 8467200, 8469000, 8470800, 
    8472600, 8474400, 8476200, 8478000, 8479800, 8481600, 8483400, 8485200, 
    8487000, 8488800, 8490600, 8492400, 8494200, 8496000, 8497800, 8499600, 
    8501400, 8503200, 8505000, 8506800, 8508600, 8510400, 8512200, 8514000, 
    8515800, 8517600, 8519400, 8521200, 8523000, 8524800, 8526600, 8528400, 
    8530200, 8532000, 8533800, 8535600, 8537400, 8539200, 8541000, 8542800, 
    8544600, 8546400, 8548200, 8550000, 8551800, 8553600, 8555400, 8557200, 
    8559000, 8560800, 8562600, 8564400, 8566200, 8568000, 8569800, 8571600, 
    8573400, 8575200, 8577000, 8578800, 8580600, 8582400, 8584200, 8586000, 
    8587800, 8589600, 8591400, 8593200, 8595000, 8596800, 8598600, 8600400, 
    8602200, 8604000, 8605800, 8607600, 8609400, 8611200, 8613000, 8614800, 
    8616600, 8618400, 8620200, 8622000, 8623800, 8625600, 8627400, 8629200, 
    8631000, 8632800, 8634600, 8636400, 8638200, 8640000, 8641800, 8643600, 
    8645400, 8647200, 8649000, 8650800, 8652600, 8654400, 8656200, 8658000, 
    8659800, 8661600, 8663400, 8665200, 8667000, 8668800, 8670600, 8672400, 
    8674200, 8676000, 8677800, 8679600, 8681400, 8683200, 8685000, 8686800, 
    8688600, 8690400, 8692200, 8694000, 8695800, 8697600, 8699400, 8701200, 
    8703000, 8704800, 8706600, 8708400, 8710200, 8712000, 8713800, 8715600, 
    8717400, 8719200, 8721000, 8722800, 8724600, 8726400, 8728200, 8730000, 
    8731800, 8733600, 8735400, 8737200, 8739000, 8740800, 8742600, 8744400, 
    8746200, 8748000, 8749800, 8751600, 8753400, 8755200, 8757000, 8758800, 
    8760600, 8762400, 8764200, 8766000, 8767800, 8769600, 8771400, 8773200, 
    8775000, 8776800, 8778600, 8780400, 8782200, 8784000, 8785800, 8787600, 
    8789400, 8791200, 8793000, 8794800, 8796600, 8798400, 8800200, 8802000, 
    8803800, 8805600, 8807400, 8809200, 8811000, 8812800, 8814600, 8816400, 
    8818200, 8820000, 8821800, 8823600, 8825400, 8827200, 8829000, 8830800, 
    8832600, 8834400, 8836200, 8838000, 8839800, 8841600, 8843400, 8845200, 
    8847000, 8848800, 8850600, 8852400, 8854200, 8856000, 8857800, 8859600, 
    8861400, 8863200, 8865000, 8866800, 8868600, 8870400, 8872200, 8874000, 
    8875800, 8877600, 8879400, 8881200, 8883000, 8884800, 8886600, 8888400, 
    8890200, 8892000, 8893800, 8895600, 8897400, 8899200, 8901000, 8902800, 
    8904600, 8906400, 8908200, 8910000, 8911800, 8913600, 8915400, 8917200, 
    8919000, 8920800, 8922600, 8924400, 8926200, 8928000, 8929800, 8931600, 
    8933400, 8935200, 8937000, 8938800, 8940600, 8942400, 8944200, 8946000, 
    8947800, 8949600, 8951400, 8953200, 8955000, 8956800, 8958600, 8960400, 
    8962200, 8964000, 8965800, 8967600, 8969400, 8971200, 8973000, 8974800, 
    8976600, 8978400, 8980200, 8982000, 8983800, 8985600, 8987400, 8989200, 
    8991000, 8992800, 8994600, 8996400, 8998200, 9000000, 9001800, 9003600, 
    9005400, 9007200, 9009000, 9010800, 9012600, 9014400, 9016200, 9018000, 
    9019800, 9021600, 9023400, 9025200, 9027000, 9028800, 9030600, 9032400, 
    9034200, 9036000, 9037800, 9039600, 9041400, 9043200, 9045000, 9046800, 
    9048600, 9050400, 9052200, 9054000, 9055800, 9057600, 9059400, 9061200, 
    9063000, 9064800, 9066600, 9068400, 9070200, 9072000, 9073800, 9075600, 
    9077400, 9079200, 9081000, 9082800, 9084600, 9086400, 9088200, 9090000, 
    9091800, 9093600, 9095400, 9097200, 9099000, 9100800, 9102600, 9104400, 
    9106200, 9108000, 9109800, 9111600, 9113400, 9115200, 9117000, 9118800, 
    9120600, 9122400, 9124200, 9126000, 9127800, 9129600, 9131400, 9133200, 
    9135000, 9136800, 9138600, 9140400, 9142200, 9144000, 9145800, 9147600, 
    9149400, 9151200, 9153000, 9154800, 9156600, 9158400, 9160200, 9162000, 
    9163800, 9165600, 9167400, 9169200, 9171000, 9172800, 9174600, 9176400, 
    9178200, 9180000, 9181800, 9183600, 9185400, 9187200, 9189000, 9190800, 
    9192600, 9194400, 9196200, 9198000, 9199800, 9201600, 9203400, 9205200, 
    9207000, 9208800, 9210600, 9212400, 9214200, 9216000, 9217800, 9219600, 
    9221400, 9223200, 9225000, 9226800, 9228600, 9230400, 9232200, 9234000, 
    9235800, 9237600, 9239400, 9241200, 9243000, 9244800, 9246600, 9248400, 
    9250200, 9252000, 9253800, 9255600, 9257400, 9259200, 9261000, 9262800, 
    9264600, 9266400, 9268200, 9270000, 9271800, 9273600, 9275400, 9277200, 
    9279000, 9280800, 9282600, 9284400, 9286200, 9288000, 9289800, 9291600, 
    9293400, 9295200, 9297000, 9298800, 9300600, 9302400, 9304200, 9306000, 
    9307800, 9309600, 9311400, 9313200, 9315000, 9316800, 9318600, 9320400, 
    9322200, 9324000, 9325800, 9327600, 9329400, 9331200, 9333000, 9334800, 
    9336600, 9338400, 9340200, 9342000, 9343800, 9345600, 9347400, 9349200, 
    9351000, 9352800, 9354600, 9356400, 9358200, 9360000, 9361800, 9363600, 
    9365400, 9367200, 9369000, 9370800, 9372600, 9374400, 9376200, 9378000, 
    9379800, 9381600, 9383400, 9385200, 9387000, 9388800, 9390600, 9392400, 
    9394200, 9396000, 9397800, 9399600, 9401400, 9403200, 9405000, 9406800, 
    9408600, 9410400, 9412200, 9414000, 9415800, 9417600, 9419400, 9421200, 
    9423000, 9424800, 9426600, 9428400, 9430200, 9432000, 9433800, 9435600, 
    9437400, 9439200, 9441000, 9442800, 9444600, 9446400, 9448200, 9450000, 
    9451800, 9453600, 9455400, 9457200, 9459000, 9460800, 9462600, 9464400, 
    9466200, 9468000, 9469800, 9471600, 9473400, 9475200, 9477000, 9478800, 
    9480600, 9482400, 9484200, 9486000, 9487800, 9489600, 9491400, 9493200, 
    9495000, 9496800, 9498600, 9500400, 9502200, 9504000, 9505800, 9507600, 
    9509400, 9511200, 9513000, 9514800, 9516600, 9518400, 9520200, 9522000, 
    9523800, 9525600, 9527400, 9529200, 9531000, 9532800, 9534600, 9536400, 
    9538200, 9540000, 9541800, 9543600, 9545400, 9547200, 9549000, 9550800, 
    9552600, 9554400, 9556200, 9558000, 9559800, 9561600, 9563400, 9565200, 
    9567000, 9568800, 9570600, 9572400, 9574200, 9576000, 9577800, 9579600, 
    9581400, 9583200, 9585000, 9586800, 9588600, 9590400, 9592200, 9594000, 
    9595800, 9597600, 9599400, 9601200, 9603000, 9604800, 9606600, 9608400, 
    9610200, 9612000, 9613800, 9615600, 9617400, 9619200, 9621000, 9622800, 
    9624600, 9626400, 9628200, 9630000, 9631800, 9633600, 9635400, 9637200, 
    9639000, 9640800, 9642600, 9644400, 9646200, 9648000, 9649800, 9651600, 
    9653400, 9655200, 9657000, 9658800, 9660600, 9662400, 9664200, 9666000, 
    9667800, 9669600, 9671400, 9673200, 9675000, 9676800, 9678600, 9680400, 
    9682200, 9684000, 9685800, 9687600, 9689400, 9691200, 9693000, 9694800, 
    9696600, 9698400, 9700200, 9702000, 9703800, 9705600, 9707400, 9709200, 
    9711000, 9712800, 9714600, 9716400, 9718200, 9720000, 9721800, 9723600, 
    9725400, 9727200, 9729000, 9730800, 9732600, 9734400, 9736200, 9738000, 
    9739800, 9741600, 9743400, 9745200, 9747000, 9748800, 9750600, 9752400, 
    9754200, 9756000, 9757800, 9759600, 9761400, 9763200, 9765000, 9766800, 
    9768600, 9770400, 9772200, 9774000, 9775800, 9777600, 9779400, 9781200, 
    9783000, 9784800, 9786600, 9788400, 9790200, 9792000, 9793800, 9795600, 
    9797400, 9799200, 9801000, 9802800, 9804600, 9806400, 9808200, 9810000, 
    9811800, 9813600, 9815400, 9817200, 9819000, 9820800, 9822600, 9824400, 
    9826200, 9828000, 9829800, 9831600, 9833400, 9835200, 9837000, 9838800, 
    9840600, 9842400, 9844200, 9846000, 9847800, 9849600, 9851400, 9853200, 
    9855000, 9856800, 9858600, 9860400, 9862200, 9864000, 9865800, 9867600, 
    9869400, 9871200, 9873000, 9874800, 9876600, 9878400, 9880200, 9882000, 
    9883800, 9885600, 9887400, 9889200, 9891000, 9892800, 9894600, 9896400, 
    9898200, 9900000, 9901800, 9903600, 9905400, 9907200, 9909000, 9910800, 
    9912600, 9914400, 9916200, 9918000, 9919800, 9921600, 9923400, 9925200, 
    9927000, 9928800, 9930600, 9932400, 9934200, 9936000, 9937800, 9939600, 
    9941400, 9943200, 9945000, 9946800, 9948600, 9950400, 9952200, 9954000, 
    9955800, 9957600, 9959400, 9961200, 9963000, 9964800, 9966600, 9968400, 
    9970200, 9972000, 9973800, 9975600, 9977400, 9979200, 9981000, 9982800, 
    9984600, 9986400, 9988200, 9990000, 9991800, 9993600, 9995400, 9997200, 
    9999000, 10000800, 10002600, 10004400, 10006200, 10008000, 10009800, 
    10011600, 10013400, 10015200, 10017000, 10018800, 10020600, 10022400, 
    10024200, 10026000, 10027800, 10029600, 10031400, 10033200, 10035000, 
    10036800, 10038600, 10040400, 10042200, 10044000, 10045800, 10047600, 
    10049400, 10051200, 10053000, 10054800, 10056600, 10058400, 10060200, 
    10062000, 10063800, 10065600, 10067400, 10069200, 10071000, 10072800, 
    10074600, 10076400, 10078200, 10080000, 10081800, 10083600, 10085400, 
    10087200, 10089000, 10090800, 10092600, 10094400, 10096200, 10098000, 
    10099800, 10101600, 10103400, 10105200, 10107000, 10108800, 10110600, 
    10112400, 10114200, 10116000, 10117800, 10119600, 10121400, 10123200, 
    10125000, 10126800, 10128600, 10130400, 10132200, 10134000, 10135800, 
    10137600, 10139400, 10141200, 10143000, 10144800, 10146600, 10148400, 
    10150200, 10152000, 10153800, 10155600, 10157400, 10159200, 10161000, 
    10162800, 10164600, 10166400, 10168200, 10170000, 10171800, 10173600, 
    10175400, 10177200, 10179000, 10180800, 10182600, 10184400, 10186200, 
    10188000, 10189800, 10191600, 10193400, 10195200, 10197000, 10198800, 
    10200600, 10202400, 10204200, 10206000, 10207800, 10209600, 10211400, 
    10213200, 10215000, 10216800, 10218600, 10220400, 10222200, 10224000, 
    10225800, 10227600, 10229400, 10231200, 10233000, 10234800, 10236600, 
    10238400, 10240200, 10242000, 10243800, 10245600, 10247400, 10249200, 
    10251000, 10252800, 10254600, 10256400, 10258200, 10260000, 10261800, 
    10263600, 10265400, 10267200, 10269000, 10270800, 10272600, 10274400, 
    10276200, 10278000, 10279800, 10281600, 10283400, 10285200, 10287000, 
    10288800, 10290600, 10292400, 10294200, 10296000, 10297800, 10299600, 
    10301400, 10303200, 10305000, 10306800, 10308600, 10310400, 10312200, 
    10314000, 10315800, 10317600, 10319400, 10321200, 10323000, 10324800, 
    10326600, 10328400, 10330200, 10332000, 10333800, 10335600, 10337400, 
    10339200, 10341000, 10342800, 10344600, 10346400, 10348200, 10350000, 
    10351800, 10353600, 10355400, 10357200, 10359000, 10360800, 10362600, 
    10364400, 10366200, 10368000, 10369800, 10371600, 10373400, 10375200, 
    10377000, 10378800, 10380600, 10382400, 10384200, 10386000, 10387800, 
    10389600, 10391400, 10393200, 10395000, 10396800, 10398600, 10400400, 
    10402200, 10404000, 10405800, 10407600, 10409400, 10411200, 10413000, 
    10414800, 10416600, 10418400, 10420200, 10422000, 10423800, 10425600, 
    10427400, 10429200, 10431000, 10432800, 10434600, 10436400, 10438200, 
    10440000, 10441800, 10443600, 10445400, 10447200, 10449000, 10450800, 
    10452600, 10454400, 10456200, 10458000, 10459800, 10461600, 10463400, 
    10465200, 10467000, 10468800, 10470600, 10472400, 10474200, 10476000, 
    10477800, 10479600, 10481400, 10483200, 10485000, 10486800, 10488600, 
    10490400, 10492200, 10494000, 10495800, 10497600, 10499400, 10501200, 
    10503000, 10504800, 10506600, 10508400, 10510200, 10512000, 10513800, 
    10515600, 10517400, 10519200, 10521000, 10522800, 10524600, 10526400, 
    10528200, 10530000, 10531800, 10533600, 10535400, 10537200, 10539000, 
    10540800, 10542600, 10544400, 10546200, 10548000, 10549800, 10551600, 
    10553400, 10555200, 10557000, 10558800, 10560600, 10562400, 10564200, 
    10566000, 10567800, 10569600, 10571400, 10573200, 10575000, 10576800, 
    10578600, 10580400, 10582200, 10584000, 10585800, 10587600, 10589400, 
    10591200, 10593000, 10594800, 10596600, 10598400, 10600200, 10602000, 
    10603800, 10605600, 10607400, 10609200, 10611000, 10612800, 10614600, 
    10616400, 10618200, 10620000, 10621800, 10623600, 10625400, 10627200, 
    10629000, 10630800, 10632600, 10634400, 10636200, 10638000, 10639800, 
    10641600, 10643400, 10645200, 10647000, 10648800, 10650600, 10652400, 
    10654200, 10656000, 10657800, 10659600, 10661400, 10663200, 10665000, 
    10666800, 10668600, 10670400, 10672200, 10674000, 10675800, 10677600, 
    10679400, 10681200, 10683000, 10684800, 10686600, 10688400, 10690200, 
    10692000, 10693800, 10695600, 10697400, 10699200, 10701000, 10702800, 
    10704600, 10706400, 10708200, 10710000, 10711800, 10713600, 10715400, 
    10717200, 10719000, 10720800, 10722600, 10724400, 10726200, 10728000, 
    10729800, 10731600, 10733400, 10735200, 10737000, 10738800, 10740600, 
    10742400, 10744200, 10746000, 10747800, 10749600, 10751400, 10753200, 
    10755000, 10756800, 10758600, 10760400, 10762200, 10764000, 10765800, 
    10767600, 10769400, 10771200, 10773000, 10774800, 10776600, 10778400, 
    10780200, 10782000, 10783800, 10785600, 10787400, 10789200, 10791000, 
    10792800, 10794600, 10796400, 10798200, 10800000, 10801800, 10803600, 
    10805400, 10807200, 10809000, 10810800, 10812600, 10814400, 10816200, 
    10818000, 10819800, 10821600, 10823400, 10825200, 10827000, 10828800, 
    10830600, 10832400, 10834200, 10836000, 10837800, 10839600, 10841400, 
    10843200, 10845000, 10846800, 10848600, 10850400, 10852200, 10854000, 
    10855800, 10857600, 10859400, 10861200, 10863000, 10864800, 10866600, 
    10868400, 10870200, 10872000, 10873800, 10875600, 10877400, 10879200, 
    10881000, 10882800, 10884600, 10886400, 10888200, 10890000, 10891800, 
    10893600, 10895400, 10897200, 10899000, 10900800, 10902600, 10904400, 
    10906200, 10908000, 10909800, 10911600, 10913400, 10915200, 10917000, 
    10918800, 10920600, 10922400, 10924200, 10926000, 10927800, 10929600, 
    10931400, 10933200, 10935000, 10936800, 10938600, 10940400, 10942200, 
    10944000, 10945800, 10947600, 10949400, 10951200, 10953000, 10954800, 
    10956600, 10958400, 10960200, 10962000, 10963800, 10965600, 10967400, 
    10969200, 10971000, 10972800, 10974600, 10976400, 10978200, 10980000, 
    10981800, 10983600, 10985400, 10987200, 10989000, 10990800, 10992600, 
    10994400, 10996200, 10998000, 10999800, 11001600, 11003400, 11005200, 
    11007000, 11008800, 11010600, 11012400, 11014200, 11016000, 11017800, 
    11019600, 11021400, 11023200, 11025000, 11026800, 11028600, 11030400, 
    11032200, 11034000, 11035800, 11037600, 11039400, 11041200, 11043000, 
    11044800, 11046600, 11048400, 11050200, 11052000, 11053800, 11055600, 
    11057400, 11059200, 11061000, 11062800, 11064600, 11066400, 11068200, 
    11070000, 11071800, 11073600, 11075400, 11077200, 11079000, 11080800, 
    11082600, 11084400, 11086200, 11088000, 11089800, 11091600, 11093400, 
    11095200, 11097000, 11098800, 11100600, 11102400, 11104200, 11106000, 
    11107800, 11109600, 11111400, 11113200, 11115000, 11116800, 11118600, 
    11120400, 11122200, 11124000, 11125800, 11127600, 11129400, 11131200, 
    11133000, 11134800, 11136600, 11138400, 11140200, 11142000, 11143800, 
    11145600, 11147400, 11149200, 11151000, 11152800, 11154600, 11156400, 
    11158200, 11160000, 11161800, 11163600, 11165400, 11167200, 11169000, 
    11170800, 11172600, 11174400, 11176200, 11178000, 11179800, 11181600, 
    11183400, 11185200, 11187000, 11188800, 11190600, 11192400, 11194200, 
    11196000, 11197800, 11199600, 11201400, 11203200, 11205000, 11206800, 
    11208600, 11210400, 11212200, 11214000, 11215800, 11217600, 11219400, 
    11221200, 11223000, 11224800, 11226600, 11228400, 11230200, 11232000, 
    11233800, 11235600, 11237400, 11239200, 11241000, 11242800, 11244600, 
    11246400, 11248200, 11250000, 11251800, 11253600, 11255400, 11257200, 
    11259000, 11260800, 11262600, 11264400, 11266200, 11268000, 11269800, 
    11271600, 11273400, 11275200, 11277000, 11278800, 11280600, 11282400, 
    11284200, 11286000, 11287800, 11289600, 11291400, 11293200, 11295000, 
    11296800, 11298600, 11300400, 11302200, 11304000, 11305800, 11307600, 
    11309400, 11311200, 11313000, 11314800, 11316600, 11318400, 11320200, 
    11322000, 11323800, 11325600, 11327400, 11329200, 11331000, 11332800, 
    11334600, 11336400, 11338200, 11340000, 11341800, 11343600, 11345400, 
    11347200, 11349000, 11350800, 11352600, 11354400, 11356200, 11358000, 
    11359800, 11361600, 11363400, 11365200, 11367000, 11368800, 11370600, 
    11372400, 11374200, 11376000, 11377800, 11379600, 11381400, 11383200, 
    11385000, 11386800, 11388600, 11390400, 11392200, 11394000, 11395800, 
    11397600, 11399400, 11401200, 11403000, 11404800, 11406600, 11408400, 
    11410200, 11412000, 11413800, 11415600, 11417400, 11419200, 11421000, 
    11422800, 11424600, 11426400, 11428200, 11430000, 11431800, 11433600, 
    11435400, 11437200, 11439000, 11440800, 11442600, 11444400, 11446200, 
    11448000, 11449800, 11451600, 11453400, 11455200, 11457000, 11458800, 
    11460600, 11462400, 11464200, 11466000, 11467800, 11469600, 11471400, 
    11473200, 11475000, 11476800, 11478600, 11480400, 11482200, 11484000, 
    11485800, 11487600, 11489400, 11491200, 11493000, 11494800, 11496600, 
    11498400, 11500200, 11502000, 11503800, 11505600, 11507400, 11509200, 
    11511000, 11512800, 11514600, 11516400, 11518200, 11520000, 11521800, 
    11523600, 11525400, 11527200, 11529000, 11530800, 11532600, 11534400, 
    11536200, 11538000, 11539800, 11541600, 11543400, 11545200, 11547000, 
    11548800, 11550600, 11552400, 11554200, 11556000, 11557800, 11559600, 
    11561400, 11563200, 11565000, 11566800, 11568600, 11570400, 11572200, 
    11574000, 11575800, 11577600, 11579400, 11581200, 11583000, 11584800, 
    11586600, 11588400, 11590200, 11592000, 11593800, 11595600, 11597400, 
    11599200, 11601000, 11602800, 11604600, 11606400, 11608200, 11610000, 
    11611800, 11613600, 11615400, 11617200, 11619000, 11620800, 11622600, 
    11624400, 11626200, 11628000, 11629800, 11631600, 11633400, 11635200, 
    11637000, 11638800, 11640600, 11642400, 11644200, 11646000, 11647800, 
    11649600, 11651400, 11653200, 11655000, 11656800, 11658600, 11660400, 
    11662200, 11664000, 11665800, 11667600, 11669400, 11671200, 11673000, 
    11674800, 11676600, 11678400, 11680200, 11682000, 11683800, 11685600, 
    11687400, 11689200, 11691000, 11692800, 11694600, 11696400, 11698200, 
    11700000, 11701800, 11703600, 11705400, 11707200, 11709000, 11710800, 
    11712600, 11714400, 11716200, 11718000, 11719800, 11721600, 11723400, 
    11725200, 11727000, 11728800, 11730600, 11732400, 11734200, 11736000, 
    11737800, 11739600, 11741400, 11743200, 11745000, 11746800, 11748600, 
    11750400, 11752200, 11754000, 11755800, 11757600, 11759400, 11761200, 
    11763000, 11764800, 11766600, 11768400, 11770200, 11772000, 11773800, 
    11775600, 11777400, 11779200, 11781000, 11782800, 11784600, 11786400, 
    11788200, 11790000, 11791800, 11793600, 11795400, 11797200, 11799000, 
    11800800, 11802600, 11804400, 11806200, 11808000, 11809800, 11811600, 
    11813400, 11815200, 11817000, 11818800, 11820600, 11822400, 11824200, 
    11826000, 11827800, 11829600, 11831400, 11833200, 11835000, 11836800, 
    11838600, 11840400, 11842200, 11844000, 11845800, 11847600, 11849400, 
    11851200, 11853000, 11854800, 11856600, 11858400, 11860200, 11862000, 
    11863800, 11865600, 11867400, 11869200, 11871000, 11872800, 11874600, 
    11876400, 11878200, 11880000, 11881800, 11883600, 11885400, 11887200, 
    11889000, 11890800, 11892600, 11894400, 11896200, 11898000, 11899800, 
    11901600, 11903400, 11905200, 11907000, 11908800, 11910600, 11912400, 
    11914200, 11916000, 11917800, 11919600, 11921400, 11923200, 11925000, 
    11926800, 11928600, 11930400, 11932200, 11934000, 11935800, 11937600, 
    11939400, 11941200, 11943000, 11944800, 11946600, 11948400, 11950200, 
    11952000, 11953800, 11955600, 11957400, 11959200, 11961000, 11962800, 
    11964600, 11966400, 11968200, 11970000, 11971800, 11973600, 11975400, 
    11977200, 11979000, 11980800, 11982600, 11984400, 11986200, 11988000, 
    11989800, 11991600, 11993400, 11995200, 11997000, 11998800, 12000600, 
    12002400, 12004200, 12006000, 12007800, 12009600, 12011400, 12013200, 
    12015000, 12016800, 12018600, 12020400, 12022200, 12024000, 12025800, 
    12027600, 12029400, 12031200, 12033000, 12034800, 12036600, 12038400, 
    12040200, 12042000, 12043800, 12045600, 12047400, 12049200, 12051000, 
    12052800, 12054600, 12056400, 12058200, 12060000, 12061800, 12063600, 
    12065400, 12067200, 12069000, 12070800, 12072600, 12074400, 12076200, 
    12078000, 12079800, 12081600, 12083400, 12085200, 12087000, 12088800, 
    12090600, 12092400, 12094200, 12096000, 12097800, 12099600, 12101400, 
    12103200, 12105000, 12106800, 12108600, 12110400, 12112200, 12114000, 
    12115800, 12117600, 12119400, 12121200, 12123000, 12124800, 12126600, 
    12128400, 12130200, 12132000, 12133800, 12135600, 12137400, 12139200, 
    12141000, 12142800, 12144600, 12146400, 12148200, 12150000, 12151800, 
    12153600, 12155400, 12157200, 12159000, 12160800, 12162600, 12164400, 
    12166200, 12168000, 12169800, 12171600, 12173400, 12175200, 12177000, 
    12178800, 12180600, 12182400, 12184200, 12186000, 12187800, 12189600, 
    12191400, 12193200, 12195000, 12196800, 12198600, 12200400, 12202200, 
    12204000, 12205800, 12207600, 12209400, 12211200, 12213000, 12214800, 
    12216600, 12218400, 12220200, 12222000, 12223800, 12225600, 12227400, 
    12229200, 12231000, 12232800, 12234600, 12236400, 12238200, 12240000, 
    12241800, 12243600, 12245400, 12247200, 12249000, 12250800, 12252600, 
    12254400, 12256200, 12258000, 12259800, 12261600, 12263400, 12265200, 
    12267000, 12268800, 12270600, 12272400, 12274200, 12276000, 12277800, 
    12279600, 12281400, 12283200, 12285000, 12286800, 12288600, 12290400, 
    12292200, 12294000, 12295800, 12297600, 12299400, 12301200, 12303000, 
    12304800, 12306600, 12308400, 12310200, 12312000, 12313800, 12315600, 
    12317400, 12319200, 12321000, 12322800, 12324600, 12326400, 12328200, 
    12330000, 12331800, 12333600, 12335400, 12337200, 12339000, 12340800, 
    12342600, 12344400, 12346200, 12348000, 12349800, 12351600, 12353400, 
    12355200, 12357000, 12358800, 12360600, 12362400, 12364200, 12366000, 
    12367800, 12369600, 12371400, 12373200, 12375000, 12376800, 12378600, 
    12380400, 12382200, 12384000, 12385800, 12387600, 12389400, 12391200, 
    12393000, 12394800, 12396600, 12398400, 12400200, 12402000, 12403800, 
    12405600, 12407400, 12409200, 12411000, 12412800, 12414600, 12416400, 
    12418200, 12420000, 12421800, 12423600, 12425400, 12427200, 12429000, 
    12430800, 12432600, 12434400, 12436200, 12438000, 12439800, 12441600, 
    12443400, 12445200, 12447000, 12448800, 12450600, 12452400, 12454200, 
    12456000, 12457800, 12459600, 12461400, 12463200, 12465000, 12466800, 
    12468600, 12470400, 12472200, 12474000, 12475800, 12477600, 12479400, 
    12481200, 12483000, 12484800, 12486600, 12488400, 12490200, 12492000, 
    12493800, 12495600, 12497400, 12499200, 12501000, 12502800, 12504600, 
    12506400, 12508200, 12510000, 12511800, 12513600, 12515400, 12517200, 
    12519000, 12520800, 12522600, 12524400, 12526200, 12528000, 12529800, 
    12531600, 12533400, 12535200, 12537000, 12538800, 12540600, 12542400, 
    12544200, 12546000, 12547800, 12549600, 12551400, 12553200, 12555000, 
    12556800, 12558600, 12560400, 12562200, 12564000, 12565800, 12567600, 
    12569400, 12571200, 12573000, 12574800, 12576600, 12578400, 12580200, 
    12582000, 12583800, 12585600, 12587400, 12589200, 12591000, 12592800, 
    12594600, 12596400, 12598200, 12600000, 12601800, 12603600, 12605400, 
    12607200, 12609000, 12610800, 12612600, 12614400, 12616200, 12618000, 
    12619800, 12621600, 12623400, 12625200, 12627000, 12628800, 12630600, 
    12632400, 12634200, 12636000, 12637800, 12639600, 12641400, 12643200, 
    12645000, 12646800, 12648600, 12650400, 12652200, 12654000, 12655800, 
    12657600, 12659400, 12661200, 12663000, 12664800, 12666600, 12668400, 
    12670200, 12672000, 12673800, 12675600, 12677400, 12679200, 12681000, 
    12682800, 12684600, 12686400, 12688200, 12690000, 12691800, 12693600, 
    12695400, 12697200, 12699000, 12700800, 12702600, 12704400, 12706200, 
    12708000, 12709800, 12711600, 12713400, 12715200, 12717000, 12718800, 
    12720600, 12722400, 12724200, 12726000, 12727800, 12729600, 12731400, 
    12733200, 12735000, 12736800, 12738600, 12740400, 12742200, 12744000, 
    12745800, 12747600, 12749400, 12751200, 12753000, 12754800, 12756600, 
    12758400, 12760200, 12762000, 12763800, 12765600, 12767400, 12769200, 
    12771000, 12772800, 12774600, 12776400, 12778200, 12780000, 12781800, 
    12783600, 12785400, 12787200, 12789000, 12790800, 12792600, 12794400, 
    12796200, 12798000, 12799800, 12801600, 12803400, 12805200, 12807000, 
    12808800, 12810600, 12812400, 12814200, 12816000, 12817800, 12819600, 
    12821400, 12823200, 12825000, 12826800, 12828600, 12830400, 12832200, 
    12834000, 12835800, 12837600, 12839400, 12841200, 12843000, 12844800, 
    12846600, 12848400, 12850200, 12852000, 12853800, 12855600, 12857400, 
    12859200, 12861000, 12862800, 12864600, 12866400, 12868200, 12870000, 
    12871800, 12873600, 12875400, 12877200, 12879000, 12880800, 12882600, 
    12884400, 12886200, 12888000, 12889800, 12891600, 12893400, 12895200, 
    12897000, 12898800, 12900600, 12902400, 12904200, 12906000, 12907800, 
    12909600, 12911400, 12913200, 12915000, 12916800, 12918600, 12920400, 
    12922200, 12924000, 12925800, 12927600, 12929400, 12931200, 12933000, 
    12934800, 12936600, 12938400, 12940200, 12942000, 12943800, 12945600, 
    12947400, 12949200, 12951000, 12952800, 12954600, 12956400, 12958200, 
    12960000, 12961800, 12963600, 12965400, 12967200, 12969000, 12970800, 
    12972600, 12974400, 12976200, 12978000, 12979800, 12981600, 12983400, 
    12985200, 12987000, 12988800, 12990600, 12992400, 12994200, 12996000, 
    12997800, 12999600, 13001400, 13003200, 13005000, 13006800, 13008600, 
    13010400, 13012200, 13014000, 13015800, 13017600, 13019400, 13021200, 
    13023000, 13024800, 13026600, 13028400, 13030200, 13032000, 13033800, 
    13035600, 13037400, 13039200, 13041000, 13042800, 13044600, 13046400, 
    13048200, 13050000, 13051800, 13053600, 13055400, 13057200, 13059000, 
    13060800, 13062600, 13064400, 13066200, 13068000, 13069800, 13071600, 
    13073400, 13075200, 13077000, 13078800, 13080600, 13082400, 13084200, 
    13086000, 13087800, 13089600, 13091400, 13093200, 13095000, 13096800, 
    13098600, 13100400, 13102200, 13104000, 13105800, 13107600, 13109400, 
    13111200, 13113000, 13114800, 13116600, 13118400, 13120200, 13122000, 
    13123800, 13125600, 13127400, 13129200, 13131000, 13132800, 13134600, 
    13136400, 13138200, 13140000, 13141800, 13143600, 13145400, 13147200, 
    13149000, 13150800, 13152600, 13154400, 13156200, 13158000, 13159800, 
    13161600, 13163400, 13165200, 13167000, 13168800, 13170600, 13172400, 
    13174200, 13176000, 13177800, 13179600, 13181400, 13183200, 13185000, 
    13186800, 13188600, 13190400, 13192200, 13194000, 13195800, 13197600, 
    13199400, 13201200, 13203000, 13204800, 13206600, 13208400, 13210200, 
    13212000, 13213800, 13215600, 13217400, 13219200, 13221000, 13222800, 
    13224600, 13226400, 13228200, 13230000, 13231800, 13233600, 13235400, 
    13237200, 13239000, 13240800, 13242600, 13244400, 13246200, 13248000, 
    13249800, 13251600, 13253400, 13255200, 13257000, 13258800, 13260600, 
    13262400, 13264200, 13266000, 13267800, 13269600, 13271400, 13273200, 
    13275000, 13276800, 13278600, 13280400, 13282200, 13284000, 13285800, 
    13287600, 13289400, 13291200, 13293000, 13294800, 13296600, 13298400, 
    13300200, 13302000, 13303800, 13305600, 13307400, 13309200, 13311000, 
    13312800, 13314600, 13316400, 13318200, 13320000, 13321800, 13323600, 
    13325400, 13327200, 13329000, 13330800, 13332600, 13334400, 13336200, 
    13338000, 13339800, 13341600, 13343400, 13345200, 13347000, 13348800, 
    13350600, 13352400, 13354200, 13356000, 13357800, 13359600, 13361400, 
    13363200, 13365000, 13366800, 13368600, 13370400, 13372200, 13374000, 
    13375800, 13377600, 13379400, 13381200, 13383000, 13384800, 13386600, 
    13388400, 13390200, 13392000, 13393800, 13395600, 13397400, 13399200, 
    13401000, 13402800, 13404600, 13406400, 13408200, 13410000, 13411800, 
    13413600, 13415400, 13417200, 13419000, 13420800, 13422600, 13424400, 
    13426200, 13428000, 13429800, 13431600, 13433400, 13435200, 13437000, 
    13438800, 13440600, 13442400, 13444200, 13446000, 13447800, 13449600, 
    13451400, 13453200, 13455000, 13456800, 13458600, 13460400, 13462200, 
    13464000, 13465800, 13467600, 13469400, 13471200, 13473000, 13474800, 
    13476600, 13478400, 13480200, 13482000, 13483800, 13485600, 13487400, 
    13489200, 13491000, 13492800, 13494600, 13496400, 13498200, 13500000, 
    13501800, 13503600, 13505400, 13507200, 13509000, 13510800, 13512600, 
    13514400, 13516200, 13518000, 13519800, 13521600, 13523400, 13525200, 
    13527000, 13528800, 13530600, 13532400, 13534200, 13536000, 13537800, 
    13539600, 13541400, 13543200, 13545000, 13546800, 13548600, 13550400, 
    13552200, 13554000, 13555800, 13557600, 13559400, 13561200, 13563000, 
    13564800, 13566600, 13568400, 13570200, 13572000, 13573800, 13575600, 
    13577400, 13579200, 13581000, 13582800, 13584600, 13586400, 13588200, 
    13590000, 13591800, 13593600, 13595400, 13597200, 13599000, 13600800, 
    13602600, 13604400, 13606200, 13608000, 13609800, 13611600, 13613400, 
    13615200, 13617000, 13618800, 13620600, 13622400, 13624200, 13626000, 
    13627800, 13629600, 13631400, 13633200, 13635000, 13636800, 13638600, 
    13640400, 13642200, 13644000, 13645800, 13647600, 13649400, 13651200, 
    13653000, 13654800, 13656600, 13658400, 13660200, 13662000, 13663800, 
    13665600, 13667400, 13669200, 13671000, 13672800, 13674600, 13676400, 
    13678200, 13680000, 13681800, 13683600, 13685400, 13687200, 13689000, 
    13690800, 13692600, 13694400, 13696200, 13698000, 13699800, 13701600, 
    13703400, 13705200, 13707000, 13708800, 13710600, 13712400, 13714200, 
    13716000, 13717800, 13719600, 13721400, 13723200, 13725000, 13726800, 
    13728600, 13730400, 13732200, 13734000, 13735800, 13737600, 13739400, 
    13741200, 13743000, 13744800, 13746600, 13748400, 13750200, 13752000, 
    13753800, 13755600, 13757400, 13759200, 13761000, 13762800, 13764600, 
    13766400, 13768200, 13770000, 13771800, 13773600, 13775400, 13777200, 
    13779000, 13780800, 13782600, 13784400, 13786200, 13788000, 13789800, 
    13791600, 13793400, 13795200, 13797000, 13798800, 13800600, 13802400, 
    13804200, 13806000, 13807800, 13809600, 13811400, 13813200, 13815000, 
    13816800, 13818600, 13820400, 13822200, 13824000, 13825800, 13827600, 
    13829400, 13831200, 13833000, 13834800, 13836600, 13838400, 13840200, 
    13842000, 13843800, 13845600, 13847400, 13849200, 13851000, 13852800, 
    13854600, 13856400, 13858200, 13860000, 13861800, 13863600, 13865400, 
    13867200, 13869000, 13870800, 13872600, 13874400, 13876200, 13878000, 
    13879800, 13881600, 13883400, 13885200, 13887000, 13888800, 13890600, 
    13892400, 13894200, 13896000, 13897800, 13899600, 13901400, 13903200, 
    13905000, 13906800, 13908600, 13910400, 13912200, 13914000, 13915800, 
    13917600, 13919400, 13921200, 13923000, 13924800, 13926600, 13928400, 
    13930200, 13932000, 13933800, 13935600, 13937400, 13939200, 13941000, 
    13942800, 13944600, 13946400, 13948200, 13950000, 13951800, 13953600, 
    13955400, 13957200, 13959000, 13960800, 13962600, 13964400, 13966200, 
    13968000, 13969800, 13971600, 13973400, 13975200, 13977000, 13978800, 
    13980600, 13982400, 13984200, 13986000, 13987800, 13989600, 13991400, 
    13993200, 13995000, 13996800, 13998600, 14000400, 14002200, 14004000, 
    14005800, 14007600, 14009400, 14011200, 14013000, 14014800, 14016600, 
    14018400, 14020200, 14022000, 14023800, 14025600, 14027400, 14029200, 
    14031000, 14032800, 14034600, 14036400, 14038200, 14040000, 14041800, 
    14043600, 14045400, 14047200, 14049000, 14050800, 14052600, 14054400, 
    14056200, 14058000, 14059800, 14061600, 14063400, 14065200, 14067000, 
    14068800, 14070600, 14072400, 14074200, 14076000, 14077800, 14079600, 
    14081400, 14083200, 14085000, 14086800, 14088600, 14090400, 14092200, 
    14094000, 14095800, 14097600, 14099400, 14101200, 14103000, 14104800, 
    14106600, 14108400, 14110200, 14112000, 14113800, 14115600, 14117400, 
    14119200, 14121000, 14122800, 14124600, 14126400, 14128200, 14130000, 
    14131800, 14133600, 14135400, 14137200, 14139000, 14140800, 14142600, 
    14144400, 14146200, 14148000, 14149800, 14151600, 14153400, 14155200, 
    14157000, 14158800, 14160600, 14162400, 14164200, 14166000, 14167800, 
    14169600, 14171400, 14173200, 14175000, 14176800, 14178600, 14180400, 
    14182200, 14184000, 14185800, 14187600, 14189400, 14191200, 14193000, 
    14194800, 14196600, 14198400, 14200200, 14202000, 14203800, 14205600, 
    14207400, 14209200, 14211000, 14212800, 14214600, 14216400, 14218200, 
    14220000, 14221800, 14223600, 14225400, 14227200, 14229000, 14230800, 
    14232600, 14234400, 14236200, 14238000, 14239800, 14241600, 14243400, 
    14245200, 14247000, 14248800, 14250600, 14252400, 14254200, 14256000, 
    14257800, 14259600, 14261400, 14263200, 14265000, 14266800, 14268600, 
    14270400, 14272200, 14274000, 14275800, 14277600, 14279400, 14281200, 
    14283000, 14284800, 14286600, 14288400, 14290200, 14292000, 14293800, 
    14295600, 14297400, 14299200, 14301000, 14302800, 14304600, 14306400, 
    14308200, 14310000, 14311800, 14313600, 14315400, 14317200, 14319000, 
    14320800, 14322600, 14324400, 14326200, 14328000, 14329800, 14331600, 
    14333400, 14335200, 14337000, 14338800, 14340600, 14342400, 14344200, 
    14346000, 14347800, 14349600, 14351400, 14353200, 14355000, 14356800, 
    14358600, 14360400, 14362200, 14364000, 14365800, 14367600, 14369400, 
    14371200, 14373000, 14374800, 14376600, 14378400, 14380200, 14382000, 
    14383800, 14385600, 14387400, 14389200, 14391000, 14392800, 14394600, 
    14396400, 14398200, 14400000, 14401800, 14403600, 14405400, 14407200, 
    14409000, 14410800, 14412600, 14414400, 14416200, 14418000, 14419800, 
    14421600, 14423400, 14425200, 14427000, 14428800, 14430600, 14432400, 
    14434200, 14436000, 14437800, 14439600, 14441400, 14443200, 14445000, 
    14446800, 14448600, 14450400, 14452200, 14454000, 14455800, 14457600, 
    14459400, 14461200, 14463000, 14464800, 14466600, 14468400, 14470200, 
    14472000, 14473800, 14475600, 14477400, 14479200, 14481000, 14482800, 
    14484600, 14486400, 14488200, 14490000, 14491800, 14493600, 14495400, 
    14497200, 14499000, 14500800, 14502600, 14504400, 14506200, 14508000, 
    14509800, 14511600, 14513400, 14515200, 14517000, 14518800, 14520600, 
    14522400, 14524200, 14526000, 14527800, 14529600, 14531400, 14533200, 
    14535000, 14536800, 14538600, 14540400, 14542200, 14544000, 14545800, 
    14547600, 14549400, 14551200, 14553000, 14554800, 14556600, 14558400, 
    14560200, 14562000, 14563800, 14565600, 14567400, 14569200, 14571000, 
    14572800, 14574600, 14576400, 14578200, 14580000, 14581800, 14583600, 
    14585400, 14587200, 14589000, 14590800, 14592600, 14594400, 14596200, 
    14598000, 14599800, 14601600, 14603400, 14605200, 14607000, 14608800, 
    14610600, 14612400, 14614200, 14616000, 14617800, 14619600, 14621400, 
    14623200, 14625000, 14626800, 14628600, 14630400, 14632200, 14634000, 
    14635800, 14637600, 14639400, 14641200, 14643000, 14644800, 14646600, 
    14648400, 14650200, 14652000, 14653800, 14655600, 14657400, 14659200, 
    14661000, 14662800, 14664600, 14666400, 14668200, 14670000, 14671800, 
    14673600, 14675400, 14677200, 14679000, 14680800, 14682600, 14684400, 
    14686200, 14688000, 14689800, 14691600, 14693400, 14695200, 14697000, 
    14698800, 14700600, 14702400, 14704200, 14706000, 14707800, 14709600, 
    14711400, 14713200, 14715000, 14716800, 14718600, 14720400, 14722200, 
    14724000, 14725800, 14727600, 14729400, 14731200, 14733000, 14734800, 
    14736600, 14738400, 14740200, 14742000, 14743800, 14745600, 14747400, 
    14749200, 14751000, 14752800, 14754600, 14756400, 14758200, 14760000, 
    14761800, 14763600, 14765400, 14767200, 14769000, 14770800, 14772600, 
    14774400, 14776200, 14778000, 14779800, 14781600, 14783400, 14785200, 
    14787000, 14788800, 14790600, 14792400, 14794200, 14796000, 14797800, 
    14799600, 14801400, 14803200, 14805000, 14806800, 14808600, 14810400, 
    14812200, 14814000, 14815800, 14817600, 14819400, 14821200, 14823000, 
    14824800, 14826600, 14828400, 14830200, 14832000, 14833800, 14835600, 
    14837400, 14839200, 14841000, 14842800, 14844600, 14846400, 14848200, 
    14850000, 14851800, 14853600, 14855400, 14857200, 14859000, 14860800, 
    14862600, 14864400, 14866200, 14868000, 14869800, 14871600, 14873400, 
    14875200, 14877000, 14878800, 14880600, 14882400, 14884200, 14886000, 
    14887800, 14889600, 14891400, 14893200, 14895000, 14896800, 14898600, 
    14900400, 14902200, 14904000, 14905800, 14907600, 14909400, 14911200, 
    14913000, 14914800, 14916600, 14918400, 14920200, 14922000, 14923800, 
    14925600, 14927400, 14929200, 14931000, 14932800, 14934600, 14936400, 
    14938200, 14940000, 14941800, 14943600, 14945400, 14947200, 14949000, 
    14950800, 14952600, 14954400, 14956200, 14958000, 14959800, 14961600, 
    14963400, 14965200, 14967000, 14968800, 14970600, 14972400, 14974200, 
    14976000, 14977800, 14979600, 14981400, 14983200, 14985000, 14986800, 
    14988600, 14990400, 14992200, 14994000, 14995800, 14997600, 14999400, 
    15001200, 15003000, 15004800, 15006600, 15008400, 15010200, 15012000, 
    15013800, 15015600, 15017400, 15019200, 15021000, 15022800, 15024600, 
    15026400, 15028200, 15030000, 15031800, 15033600, 15035400, 15037200, 
    15039000, 15040800, 15042600, 15044400, 15046200, 15048000, 15049800, 
    15051600, 15053400, 15055200, 15057000, 15058800, 15060600, 15062400, 
    15064200, 15066000, 15067800, 15069600, 15071400, 15073200, 15075000, 
    15076800, 15078600, 15080400, 15082200, 15084000, 15085800, 15087600, 
    15089400, 15091200, 15093000, 15094800, 15096600, 15098400, 15100200, 
    15102000, 15103800, 15105600, 15107400, 15109200, 15111000, 15112800, 
    15114600, 15116400, 15118200, 15120000, 15121800, 15123600, 15125400, 
    15127200, 15129000, 15130800, 15132600, 15134400, 15136200, 15138000, 
    15139800, 15141600, 15143400, 15145200, 15147000, 15148800, 15150600, 
    15152400, 15154200, 15156000, 15157800, 15159600, 15161400, 15163200, 
    15165000, 15166800, 15168600, 15170400, 15172200, 15174000, 15175800, 
    15177600, 15179400, 15181200, 15183000, 15184800, 15186600, 15188400, 
    15190200, 15192000, 15193800, 15195600, 15197400, 15199200, 15201000, 
    15202800, 15204600, 15206400, 15208200, 15210000, 15211800, 15213600, 
    15215400, 15217200, 15219000, 15220800, 15222600, 15224400, 15226200, 
    15228000, 15229800, 15231600, 15233400, 15235200, 15237000, 15238800, 
    15240600, 15242400, 15244200, 15246000, 15247800, 15249600, 15251400, 
    15253200, 15255000, 15256800, 15258600, 15260400, 15262200, 15264000, 
    15265800, 15267600, 15269400, 15271200, 15273000, 15274800, 15276600, 
    15278400, 15280200, 15282000, 15283800, 15285600, 15287400, 15289200, 
    15291000, 15292800, 15294600, 15296400, 15298200, 15300000, 15301800, 
    15303600, 15305400, 15307200, 15309000, 15310800, 15312600, 15314400, 
    15316200, 15318000, 15319800, 15321600, 15323400, 15325200, 15327000, 
    15328800, 15330600, 15332400, 15334200, 15336000, 15337800, 15339600, 
    15341400, 15343200, 15345000, 15346800, 15348600, 15350400, 15352200, 
    15354000, 15355800, 15357600, 15359400, 15361200, 15363000, 15364800, 
    15366600, 15368400, 15370200, 15372000, 15373800, 15375600, 15377400, 
    15379200, 15381000, 15382800, 15384600, 15386400, 15388200, 15390000, 
    15391800, 15393600, 15395400, 15397200, 15399000, 15400800, 15402600, 
    15404400, 15406200, 15408000, 15409800, 15411600, 15413400, 15415200, 
    15417000, 15418800, 15420600, 15422400, 15424200, 15426000, 15427800, 
    15429600, 15431400, 15433200, 15435000, 15436800, 15438600, 15440400, 
    15442200, 15444000, 15445800, 15447600, 15449400, 15451200, 15453000, 
    15454800, 15456600, 15458400, 15460200, 15462000, 15463800, 15465600, 
    15467400, 15469200, 15471000, 15472800, 15474600, 15476400, 15478200, 
    15480000, 15481800, 15483600, 15485400, 15487200, 15489000, 15490800, 
    15492600, 15494400, 15496200, 15498000, 15499800, 15501600, 15503400, 
    15505200, 15507000, 15508800, 15510600, 15512400, 15514200, 15516000, 
    15517800, 15519600, 15521400, 15523200, 15525000, 15526800, 15528600, 
    15530400, 15532200, 15534000, 15535800, 15537600, 15539400, 15541200, 
    15543000, 15544800, 15546600, 15548400, 15550200, 15552000, 15553800, 
    15555600, 15557400, 15559200, 15561000, 15562800, 15564600, 15566400, 
    15568200, 15570000, 15571800, 15573600, 15575400, 15577200, 15579000, 
    15580800, 15582600, 15584400, 15586200, 15588000, 15589800, 15591600, 
    15593400, 15595200, 15597000, 15598800, 15600600, 15602400, 15604200, 
    15606000, 15607800, 15609600, 15611400, 15613200, 15615000, 15616800, 
    15618600, 15620400, 15622200, 15624000, 15625800, 15627600, 15629400, 
    15631200, 15633000, 15634800, 15636600, 15638400, 15640200, 15642000, 
    15643800, 15645600, 15647400, 15649200, 15651000, 15652800, 15654600, 
    15656400, 15658200, 15660000, 15661800, 15663600, 15665400, 15667200, 
    15669000, 15670800, 15672600, 15674400, 15676200, 15678000, 15679800, 
    15681600, 15683400, 15685200, 15687000, 15688800, 15690600, 15692400, 
    15694200, 15696000, 15697800, 15699600, 15701400, 15703200, 15705000, 
    15706800, 15708600, 15710400, 15712200, 15714000, 15715800, 15717600, 
    15719400, 15721200, 15723000, 15724800, 15726600, 15728400, 15730200, 
    15732000, 15733800, 15735600, 15737400, 15739200, 15741000, 15742800, 
    15744600, 15746400, 15748200, 15750000, 15751800, 15753600, 15755400, 
    15757200, 15759000, 15760800, 15762600, 15764400, 15766200, 15768000, 
    15769800, 15771600, 15773400, 15775200, 15777000, 15778800, 15780600, 
    15782400, 15784200, 15786000, 15787800, 15789600, 15791400, 15793200, 
    15795000, 15796800, 15798600, 15800400, 15802200, 15804000, 15805800, 
    15807600, 15809400, 15811200, 15813000, 15814800, 15816600, 15818400, 
    15820200, 15822000, 15823800, 15825600, 15827400, 15829200, 15831000, 
    15832800, 15834600, 15836400, 15838200, 15840000, 15841800, 15843600, 
    15845400, 15847200, 15849000, 15850800, 15852600, 15854400, 15856200, 
    15858000, 15859800, 15861600, 15863400, 15865200, 15867000, 15868800, 
    15870600, 15872400, 15874200, 15876000, 15877800, 15879600, 15881400, 
    15883200, 15885000, 15886800, 15888600, 15890400, 15892200, 15894000, 
    15895800, 15897600, 15899400, 15901200, 15903000, 15904800, 15906600, 
    15908400, 15910200, 15912000, 15913800, 15915600, 15917400, 15919200, 
    15921000, 15922800, 15924600, 15926400, 15928200, 15930000, 15931800, 
    15933600, 15935400, 15937200, 15939000, 15940800, 15942600, 15944400, 
    15946200, 15948000, 15949800, 15951600, 15953400, 15955200, 15957000, 
    15958800, 15960600, 15962400, 15964200, 15966000, 15967800, 15969600, 
    15971400, 15973200, 15975000, 15976800, 15978600, 15980400, 15982200, 
    15984000, 15985800, 15987600, 15989400, 15991200, 15993000, 15994800, 
    15996600, 15998400, 16000200, 16002000, 16003800, 16005600, 16007400, 
    16009200, 16011000, 16012800, 16014600, 16016400, 16018200, 16020000, 
    16021800, 16023600, 16025400, 16027200, 16029000, 16030800, 16032600, 
    16034400, 16036200, 16038000, 16039800, 16041600, 16043400, 16045200, 
    16047000, 16048800, 16050600, 16052400, 16054200, 16056000, 16057800, 
    16059600, 16061400, 16063200, 16065000, 16066800, 16068600, 16070400, 
    16072200, 16074000, 16075800, 16077600, 16079400, 16081200, 16083000, 
    16084800, 16086600, 16088400, 16090200, 16092000, 16093800, 16095600, 
    16097400, 16099200, 16101000, 16102800, 16104600, 16106400, 16108200, 
    16110000, 16111800, 16113600, 16115400, 16117200, 16119000, 16120800, 
    16122600, 16124400, 16126200, 16128000, 16129800, 16131600, 16133400, 
    16135200, 16137000, 16138800, 16140600, 16142400, 16144200, 16146000, 
    16147800, 16149600, 16151400, 16153200, 16155000, 16156800, 16158600, 
    16160400, 16162200, 16164000, 16165800, 16167600, 16169400, 16171200, 
    16173000, 16174800, 16176600, 16178400, 16180200, 16182000, 16183800, 
    16185600, 16187400, 16189200, 16191000, 16192800, 16194600, 16196400, 
    16198200, 16200000, 16201800, 16203600, 16205400, 16207200, 16209000, 
    16210800, 16212600, 16214400, 16216200, 16218000, 16219800, 16221600, 
    16223400, 16225200, 16227000, 16228800, 16230600, 16232400, 16234200, 
    16236000, 16237800, 16239600, 16241400, 16243200, 16245000, 16246800, 
    16248600, 16250400, 16252200, 16254000, 16255800, 16257600, 16259400, 
    16261200, 16263000, 16264800, 16266600, 16268400, 16270200, 16272000, 
    16273800, 16275600, 16277400, 16279200, 16281000, 16282800, 16284600, 
    16286400, 16288200, 16290000, 16291800, 16293600, 16295400, 16297200, 
    16299000, 16300800, 16302600, 16304400, 16306200, 16308000, 16309800, 
    16311600, 16313400, 16315200, 16317000, 16318800, 16320600, 16322400, 
    16324200, 16326000, 16327800, 16329600, 16331400, 16333200, 16335000, 
    16336800, 16338600, 16340400, 16342200, 16344000, 16345800, 16347600, 
    16349400, 16351200, 16353000, 16354800, 16356600, 16358400, 16360200, 
    16362000, 16363800, 16365600, 16367400, 16369200, 16371000, 16372800, 
    16374600, 16376400, 16378200, 16380000, 16381800, 16383600, 16385400, 
    16387200, 16389000, 16390800, 16392600, 16394400, 16396200, 16398000, 
    16399800, 16401600, 16403400, 16405200, 16407000, 16408800, 16410600, 
    16412400, 16414200, 16416000, 16417800, 16419600, 16421400, 16423200, 
    16425000, 16426800, 16428600, 16430400, 16432200, 16434000, 16435800, 
    16437600, 16439400, 16441200, 16443000, 16444800, 16446600, 16448400, 
    16450200, 16452000, 16453800, 16455600, 16457400, 16459200, 16461000, 
    16462800, 16464600, 16466400, 16468200, 16470000, 16471800, 16473600, 
    16475400, 16477200, 16479000, 16480800, 16482600, 16484400, 16486200, 
    16488000, 16489800, 16491600, 16493400, 16495200, 16497000, 16498800, 
    16500600, 16502400, 16504200, 16506000, 16507800, 16509600, 16511400, 
    16513200, 16515000, 16516800, 16518600, 16520400, 16522200, 16524000, 
    16525800, 16527600, 16529400, 16531200, 16533000, 16534800, 16536600, 
    16538400, 16540200, 16542000, 16543800, 16545600, 16547400, 16549200, 
    16551000, 16552800, 16554600, 16556400, 16558200, 16560000, 16561800, 
    16563600, 16565400, 16567200, 16569000, 16570800, 16572600, 16574400, 
    16576200, 16578000, 16579800, 16581600, 16583400, 16585200, 16587000, 
    16588800, 16590600, 16592400, 16594200, 16596000, 16597800, 16599600, 
    16601400, 16603200, 16605000, 16606800, 16608600, 16610400, 16612200, 
    16614000, 16615800, 16617600, 16619400, 16621200, 16623000, 16624800, 
    16626600, 16628400, 16630200, 16632000, 16633800, 16635600, 16637400, 
    16639200, 16641000, 16642800, 16644600, 16646400, 16648200, 16650000, 
    16651800, 16653600, 16655400, 16657200, 16659000, 16660800, 16662600, 
    16664400, 16666200, 16668000, 16669800, 16671600, 16673400, 16675200, 
    16677000, 16678800, 16680600, 16682400, 16684200, 16686000, 16687800, 
    16689600, 16691400, 16693200, 16695000, 16696800, 16698600, 16700400, 
    16702200, 16704000, 16705800, 16707600, 16709400, 16711200, 16713000, 
    16714800, 16716600, 16718400, 16720200, 16722000, 16723800, 16725600, 
    16727400, 16729200, 16731000, 16732800, 16734600, 16736400, 16738200, 
    16740000, 16741800, 16743600, 16745400, 16747200, 16749000, 16750800, 
    16752600, 16754400, 16756200, 16758000, 16759800, 16761600, 16763400, 
    16765200, 16767000, 16768800, 16770600, 16772400, 16774200, 16776000, 
    16777800, 16779600, 16781400, 16783200, 16785000, 16786800, 16788600, 
    16790400, 16792200, 16794000, 16795800, 16797600, 16799400, 16801200, 
    16803000, 16804800, 16806600, 16808400, 16810200, 16812000, 16813800, 
    16815600, 16817400, 16819200, 16821000, 16822800, 16824600, 16826400, 
    16828200, 16830000, 16831800, 16833600, 16835400, 16837200, 16839000, 
    16840800, 16842600, 16844400, 16846200, 16848000, 16849800, 16851600, 
    16853400, 16855200, 16857000, 16858800, 16860600, 16862400, 16864200, 
    16866000, 16867800, 16869600, 16871400, 16873200, 16875000, 16876800, 
    16878600, 16880400, 16882200, 16884000, 16885800, 16887600, 16889400, 
    16891200, 16893000, 16894800, 16896600, 16898400, 16900200, 16902000, 
    16903800, 16905600, 16907400, 16909200, 16911000, 16912800, 16914600, 
    16916400, 16918200, 16920000, 16921800, 16923600, 16925400, 16927200, 
    16929000, 16930800, 16932600, 16934400, 16936200, 16938000, 16939800, 
    16941600, 16943400, 16945200, 16947000, 16948800, 16950600, 16952400, 
    16954200, 16956000, 16957800, 16959600, 16961400, 16963200, 16965000, 
    16966800, 16968600, 16970400, 16972200, 16974000, 16975800, 16977600, 
    16979400, 16981200, 16983000, 16984800, 16986600, 16988400, 16990200, 
    16992000, 16993800, 16995600, 16997400, 16999200, 17001000, 17002800, 
    17004600, 17006400, 17008200, 17010000, 17011800, 17013600, 17015400, 
    17017200, 17019000, 17020800, 17022600, 17024400, 17026200, 17028000, 
    17029800, 17031600, 17033400, 17035200, 17037000, 17038800, 17040600, 
    17042400, 17044200, 17046000, 17047800, 17049600, 17051400, 17053200, 
    17055000, 17056800, 17058600, 17060400, 17062200, 17064000, 17065800, 
    17067600, 17069400, 17071200, 17073000, 17074800, 17076600, 17078400, 
    17080200, 17082000, 17083800, 17085600, 17087400, 17089200, 17091000, 
    17092800, 17094600, 17096400, 17098200, 17100000, 17101800, 17103600, 
    17105400, 17107200, 17109000, 17110800, 17112600, 17114400, 17116200, 
    17118000, 17119800, 17121600, 17123400, 17125200, 17127000, 17128800, 
    17130600, 17132400, 17134200, 17136000, 17137800, 17139600, 17141400, 
    17143200, 17145000, 17146800, 17148600, 17150400, 17152200, 17154000, 
    17155800, 17157600, 17159400, 17161200, 17163000, 17164800, 17166600, 
    17168400, 17170200, 17172000, 17173800, 17175600, 17177400, 17179200, 
    17181000, 17182800, 17184600, 17186400, 17188200, 17190000, 17191800, 
    17193600, 17195400, 17197200, 17199000, 17200800, 17202600, 17204400, 
    17206200, 17208000, 17209800, 17211600, 17213400, 17215200, 17217000, 
    17218800, 17220600, 17222400, 17224200, 17226000, 17227800, 17229600, 
    17231400, 17233200, 17235000, 17236800, 17238600, 17240400, 17242200, 
    17244000, 17245800, 17247600, 17249400, 17251200, 17253000, 17254800, 
    17256600, 17258400, 17260200, 17262000, 17263800, 17265600, 17267400, 
    17269200, 17271000, 17272800, 17274600, 17276400, 17278200, 17280000, 
    17281800, 17283600, 17285400, 17287200, 17289000, 17290800, 17292600, 
    17294400, 17296200, 17298000, 17299800, 17301600, 17303400, 17305200, 
    17307000, 17308800, 17310600, 17312400, 17314200, 17316000, 17317800, 
    17319600, 17321400, 17323200, 17325000, 17326800, 17328600, 17330400, 
    17332200, 17334000, 17335800, 17337600, 17339400, 17341200, 17343000, 
    17344800, 17346600, 17348400, 17350200, 17352000, 17353800, 17355600, 
    17357400, 17359200, 17361000, 17362800, 17364600, 17366400, 17368200, 
    17370000, 17371800, 17373600, 17375400, 17377200, 17379000, 17380800, 
    17382600, 17384400, 17386200, 17388000, 17389800, 17391600, 17393400, 
    17395200, 17397000, 17398800, 17400600, 17402400, 17404200, 17406000, 
    17407800, 17409600, 17411400, 17413200, 17415000, 17416800, 17418600, 
    17420400, 17422200, 17424000, 17425800, 17427600, 17429400, 17431200, 
    17433000, 17434800, 17436600, 17438400, 17440200, 17442000, 17443800, 
    17445600, 17447400, 17449200, 17451000, 17452800, 17454600, 17456400, 
    17458200, 17460000, 17461800, 17463600, 17465400, 17467200, 17469000, 
    17470800, 17472600, 17474400, 17476200, 17478000, 17479800, 17481600, 
    17483400, 17485200, 17487000, 17488800, 17490600, 17492400, 17494200, 
    17496000, 17497800, 17499600, 17501400, 17503200, 17505000, 17506800, 
    17508600, 17510400, 17512200, 17514000, 17515800, 17517600, 17519400, 
    17521200, 17523000, 17524800, 17526600, 17528400, 17530200, 17532000, 
    17533800, 17535600, 17537400, 17539200, 17541000, 17542800, 17544600, 
    17546400, 17548200, 17550000, 17551800, 17553600, 17555400, 17557200, 
    17559000, 17560800, 17562600, 17564400, 17566200, 17568000, 17569800, 
    17571600, 17573400, 17575200, 17577000, 17578800, 17580600, 17582400, 
    17584200, 17586000, 17587800, 17589600, 17591400, 17593200, 17595000, 
    17596800, 17598600, 17600400, 17602200, 17604000, 17605800, 17607600, 
    17609400, 17611200, 17613000, 17614800, 17616600, 17618400, 17620200, 
    17622000, 17623800, 17625600, 17627400, 17629200, 17631000, 17632800, 
    17634600, 17636400, 17638200, 17640000, 17641800, 17643600, 17645400, 
    17647200, 17649000, 17650800, 17652600, 17654400, 17656200, 17658000, 
    17659800, 17661600, 17663400, 17665200, 17667000, 17668800, 17670600, 
    17672400, 17674200, 17676000, 17677800, 17679600, 17681400, 17683200, 
    17685000, 17686800, 17688600, 17690400, 17692200, 17694000, 17695800, 
    17697600, 17699400, 17701200, 17703000, 17704800, 17706600, 17708400, 
    17710200, 17712000, 17713800, 17715600, 17717400, 17719200, 17721000, 
    17722800, 17724600, 17726400, 17728200, 17730000, 17731800, 17733600, 
    17735400, 17737200, 17739000, 17740800, 17742600, 17744400, 17746200, 
    17748000, 17749800, 17751600, 17753400, 17755200, 17757000, 17758800, 
    17760600, 17762400, 17764200, 17766000, 17767800, 17769600, 17771400, 
    17773200, 17775000, 17776800, 17778600, 17780400, 17782200, 17784000, 
    17785800, 17787600, 17789400, 17791200, 17793000, 17794800, 17796600, 
    17798400, 17800200, 17802000, 17803800, 17805600, 17807400, 17809200, 
    17811000, 17812800, 17814600, 17816400, 17818200, 17820000, 17821800, 
    17823600, 17825400, 17827200, 17829000, 17830800, 17832600, 17834400, 
    17836200, 17838000, 17839800, 17841600, 17843400, 17845200, 17847000, 
    17848800, 17850600, 17852400, 17854200, 17856000, 17857800, 17859600, 
    17861400, 17863200, 17865000, 17866800, 17868600, 17870400, 17872200, 
    17874000, 17875800, 17877600, 17879400, 17881200, 17883000, 17884800, 
    17886600, 17888400, 17890200, 17892000, 17893800, 17895600, 17897400, 
    17899200, 17901000, 17902800, 17904600, 17906400, 17908200, 17910000, 
    17911800, 17913600, 17915400, 17917200, 17919000, 17920800, 17922600, 
    17924400, 17926200, 17928000, 17929800, 17931600, 17933400, 17935200, 
    17937000, 17938800, 17940600, 17942400, 17944200, 17946000, 17947800, 
    17949600, 17951400, 17953200, 17955000, 17956800, 17958600, 17960400, 
    17962200, 17964000, 17965800, 17967600, 17969400, 17971200, 17973000, 
    17974800, 17976600, 17978400, 17980200, 17982000, 17983800, 17985600, 
    17987400, 17989200, 17991000, 17992800, 17994600, 17996400, 17998200, 
    18000000, 18001800, 18003600, 18005400, 18007200, 18009000, 18010800, 
    18012600, 18014400, 18016200, 18018000, 18019800, 18021600, 18023400, 
    18025200, 18027000, 18028800, 18030600, 18032400, 18034200, 18036000, 
    18037800, 18039600, 18041400, 18043200, 18045000, 18046800, 18048600, 
    18050400, 18052200, 18054000, 18055800, 18057600, 18059400, 18061200, 
    18063000, 18064800, 18066600, 18068400, 18070200, 18072000, 18073800, 
    18075600, 18077400, 18079200, 18081000, 18082800, 18084600, 18086400, 
    18088200, 18090000, 18091800, 18093600, 18095400, 18097200, 18099000, 
    18100800, 18102600, 18104400, 18106200, 18108000, 18109800, 18111600, 
    18113400, 18115200, 18117000, 18118800, 18120600, 18122400, 18124200, 
    18126000, 18127800, 18129600, 18131400, 18133200, 18135000, 18136800, 
    18138600, 18140400, 18142200, 18144000, 18145800, 18147600, 18149400, 
    18151200, 18153000, 18154800, 18156600, 18158400, 18160200, 18162000, 
    18163800, 18165600, 18167400, 18169200, 18171000, 18172800, 18174600, 
    18176400, 18178200, 18180000, 18181800, 18183600, 18185400, 18187200, 
    18189000, 18190800, 18192600, 18194400, 18196200, 18198000, 18199800, 
    18201600, 18203400, 18205200, 18207000, 18208800, 18210600, 18212400, 
    18214200, 18216000, 18217800, 18219600, 18221400, 18223200, 18225000, 
    18226800, 18228600, 18230400, 18232200, 18234000, 18235800, 18237600, 
    18239400, 18241200, 18243000, 18244800, 18246600, 18248400, 18250200, 
    18252000, 18253800, 18255600, 18257400, 18259200, 18261000, 18262800, 
    18264600, 18266400, 18268200, 18270000, 18271800, 18273600, 18275400, 
    18277200, 18279000, 18280800, 18282600, 18284400, 18286200, 18288000, 
    18289800, 18291600, 18293400, 18295200, 18297000, 18298800, 18300600, 
    18302400, 18304200, 18306000, 18307800, 18309600, 18311400, 18313200, 
    18315000, 18316800, 18318600, 18320400, 18322200, 18324000, 18325800, 
    18327600, 18329400, 18331200, 18333000, 18334800, 18336600, 18338400, 
    18340200, 18342000, 18343800, 18345600, 18347400, 18349200, 18351000, 
    18352800, 18354600, 18356400, 18358200, 18360000, 18361800, 18363600, 
    18365400, 18367200, 18369000, 18370800, 18372600, 18374400, 18376200, 
    18378000, 18379800, 18381600, 18383400, 18385200, 18387000, 18388800, 
    18390600, 18392400, 18394200, 18396000, 18397800, 18399600, 18401400, 
    18403200, 18405000, 18406800, 18408600, 18410400, 18412200, 18414000, 
    18415800, 18417600, 18419400, 18421200, 18423000, 18424800, 18426600, 
    18428400, 18430200, 18432000, 18433800, 18435600, 18437400, 18439200, 
    18441000, 18442800, 18444600, 18446400, 18448200, 18450000, 18451800, 
    18453600, 18455400, 18457200, 18459000, 18460800, 18462600, 18464400, 
    18466200, 18468000, 18469800, 18471600, 18473400, 18475200, 18477000, 
    18478800, 18480600, 18482400, 18484200, 18486000, 18487800, 18489600, 
    18491400, 18493200, 18495000, 18496800, 18498600, 18500400, 18502200, 
    18504000, 18505800, 18507600, 18509400, 18511200, 18513000, 18514800, 
    18516600, 18518400, 18520200, 18522000, 18523800, 18525600, 18527400, 
    18529200, 18531000, 18532800, 18534600, 18536400, 18538200, 18540000, 
    18541800, 18543600, 18545400, 18547200, 18549000, 18550800, 18552600, 
    18554400, 18556200, 18558000, 18559800, 18561600, 18563400, 18565200, 
    18567000, 18568800, 18570600, 18572400, 18574200, 18576000, 18577800, 
    18579600, 18581400, 18583200, 18585000, 18586800, 18588600, 18590400, 
    18592200, 18594000, 18595800, 18597600, 18599400, 18601200, 18603000, 
    18604800, 18606600, 18608400, 18610200, 18612000, 18613800, 18615600, 
    18617400, 18619200, 18621000, 18622800, 18624600, 18626400, 18628200, 
    18630000, 18631800, 18633600, 18635400, 18637200, 18639000, 18640800, 
    18642600, 18644400, 18646200, 18648000, 18649800, 18651600, 18653400, 
    18655200, 18657000, 18658800, 18660600, 18662400, 18664200, 18666000, 
    18667800, 18669600, 18671400, 18673200, 18675000, 18676800, 18678600, 
    18680400, 18682200, 18684000, 18685800, 18687600, 18689400, 18691200, 
    18693000, 18694800, 18696600, 18698400, 18700200, 18702000, 18703800, 
    18705600, 18707400, 18709200, 18711000, 18712800, 18714600, 18716400, 
    18718200, 18720000, 18721800, 18723600, 18725400, 18727200, 18729000, 
    18730800, 18732600, 18734400, 18736200, 18738000, 18739800, 18741600, 
    18743400, 18745200, 18747000, 18748800, 18750600, 18752400, 18754200, 
    18756000, 18757800, 18759600, 18761400, 18763200, 18765000, 18766800, 
    18768600, 18770400, 18772200, 18774000, 18775800, 18777600, 18779400, 
    18781200, 18783000, 18784800, 18786600, 18788400, 18790200, 18792000, 
    18793800, 18795600, 18797400, 18799200, 18801000, 18802800, 18804600, 
    18806400, 18808200, 18810000, 18811800, 18813600, 18815400, 18817200, 
    18819000, 18820800, 18822600, 18824400, 18826200, 18828000, 18829800, 
    18831600, 18833400, 18835200, 18837000, 18838800, 18840600, 18842400, 
    18844200, 18846000, 18847800, 18849600, 18851400, 18853200, 18855000, 
    18856800, 18858600, 18860400, 18862200, 18864000, 18865800, 18867600, 
    18869400, 18871200, 18873000, 18874800, 18876600, 18878400, 18880200, 
    18882000, 18883800, 18885600, 18887400, 18889200, 18891000, 18892800, 
    18894600, 18896400, 18898200, 18900000, 18901800, 18903600, 18905400, 
    18907200, 18909000, 18910800, 18912600, 18914400, 18916200, 18918000, 
    18919800, 18921600, 18923400, 18925200, 18927000, 18928800, 18930600, 
    18932400, 18934200, 18936000, 18937800, 18939600, 18941400, 18943200, 
    18945000, 18946800, 18948600, 18950400, 18952200, 18954000, 18955800, 
    18957600, 18959400, 18961200, 18963000, 18964800, 18966600, 18968400, 
    18970200, 18972000, 18973800, 18975600, 18977400, 18979200, 18981000, 
    18982800, 18984600, 18986400, 18988200, 18990000, 18991800, 18993600, 
    18995400, 18997200, 18999000, 19000800, 19002600, 19004400, 19006200, 
    19008000, 19009800, 19011600, 19013400, 19015200, 19017000, 19018800, 
    19020600, 19022400, 19024200, 19026000, 19027800, 19029600, 19031400, 
    19033200, 19035000, 19036800, 19038600, 19040400, 19042200, 19044000, 
    19045800, 19047600, 19049400, 19051200, 19053000, 19054800, 19056600, 
    19058400, 19060200, 19062000, 19063800, 19065600, 19067400, 19069200, 
    19071000, 19072800, 19074600, 19076400, 19078200, 19080000, 19081800, 
    19083600, 19085400, 19087200, 19089000, 19090800, 19092600, 19094400, 
    19096200, 19098000, 19099800, 19101600, 19103400, 19105200, 19107000, 
    19108800, 19110600, 19112400, 19114200, 19116000, 19117800, 19119600, 
    19121400, 19123200, 19125000, 19126800, 19128600, 19130400, 19132200, 
    19134000, 19135800, 19137600, 19139400, 19141200, 19143000, 19144800, 
    19146600, 19148400, 19150200, 19152000, 19153800, 19155600, 19157400, 
    19159200, 19161000, 19162800, 19164600, 19166400, 19168200, 19170000, 
    19171800, 19173600, 19175400, 19177200, 19179000, 19180800, 19182600, 
    19184400, 19186200, 19188000, 19189800, 19191600, 19193400, 19195200, 
    19197000, 19198800, 19200600, 19202400, 19204200, 19206000, 19207800, 
    19209600, 19211400, 19213200, 19215000, 19216800, 19218600, 19220400, 
    19222200, 19224000, 19225800, 19227600, 19229400, 19231200, 19233000, 
    19234800, 19236600, 19238400, 19240200, 19242000, 19243800, 19245600, 
    19247400, 19249200, 19251000, 19252800, 19254600, 19256400, 19258200, 
    19260000, 19261800, 19263600, 19265400, 19267200, 19269000, 19270800, 
    19272600, 19274400, 19276200, 19278000, 19279800, 19281600, 19283400, 
    19285200, 19287000, 19288800, 19290600, 19292400, 19294200, 19296000, 
    19297800, 19299600, 19301400, 19303200, 19305000, 19306800, 19308600, 
    19310400, 19312200, 19314000, 19315800, 19317600, 19319400, 19321200, 
    19323000, 19324800, 19326600, 19328400, 19330200, 19332000, 19333800, 
    19335600, 19337400, 19339200, 19341000, 19342800, 19344600, 19346400, 
    19348200, 19350000, 19351800, 19353600, 19355400, 19357200, 19359000, 
    19360800, 19362600, 19364400, 19366200, 19368000, 19369800, 19371600, 
    19373400, 19375200, 19377000, 19378800, 19380600, 19382400, 19384200, 
    19386000, 19387800, 19389600, 19391400, 19393200, 19395000, 19396800, 
    19398600, 19400400, 19402200, 19404000, 19405800, 19407600, 19409400, 
    19411200, 19413000, 19414800, 19416600, 19418400, 19420200, 19422000, 
    19423800, 19425600, 19427400, 19429200, 19431000, 19432800, 19434600, 
    19436400, 19438200, 19440000, 19441800, 19443600, 19445400, 19447200, 
    19449000, 19450800, 19452600, 19454400, 19456200, 19458000, 19459800, 
    19461600, 19463400, 19465200, 19467000, 19468800, 19470600, 19472400, 
    19474200, 19476000, 19477800, 19479600, 19481400, 19483200, 19485000, 
    19486800, 19488600, 19490400, 19492200, 19494000, 19495800, 19497600, 
    19499400, 19501200, 19503000, 19504800, 19506600, 19508400, 19510200, 
    19512000, 19513800, 19515600, 19517400, 19519200, 19521000, 19522800, 
    19524600, 19526400, 19528200, 19530000, 19531800, 19533600, 19535400, 
    19537200, 19539000, 19540800, 19542600, 19544400, 19546200, 19548000, 
    19549800, 19551600, 19553400, 19555200, 19557000, 19558800, 19560600, 
    19562400, 19564200, 19566000, 19567800, 19569600, 19571400, 19573200, 
    19575000, 19576800, 19578600, 19580400, 19582200, 19584000, 19585800, 
    19587600, 19589400, 19591200, 19593000, 19594800, 19596600, 19598400, 
    19600200, 19602000, 19603800, 19605600, 19607400, 19609200, 19611000, 
    19612800, 19614600, 19616400, 19618200, 19620000, 19621800, 19623600, 
    19625400, 19627200, 19629000, 19630800, 19632600, 19634400, 19636200, 
    19638000, 19639800, 19641600, 19643400, 19645200, 19647000, 19648800, 
    19650600, 19652400, 19654200, 19656000, 19657800, 19659600, 19661400, 
    19663200, 19665000, 19666800, 19668600, 19670400, 19672200, 19674000, 
    19675800, 19677600, 19679400, 19681200, 19683000, 19684800, 19686600, 
    19688400, 19690200, 19692000, 19693800, 19695600, 19697400, 19699200, 
    19701000, 19702800, 19704600, 19706400, 19708200, 19710000, 19711800, 
    19713600, 19715400, 19717200, 19719000, 19720800, 19722600, 19724400, 
    19726200, 19728000, 19729800, 19731600, 19733400, 19735200, 19737000, 
    19738800, 19740600, 19742400, 19744200, 19746000, 19747800, 19749600, 
    19751400, 19753200, 19755000, 19756800, 19758600, 19760400, 19762200, 
    19764000, 19765800, 19767600, 19769400, 19771200, 19773000, 19774800, 
    19776600, 19778400, 19780200, 19782000, 19783800, 19785600, 19787400, 
    19789200, 19791000, 19792800, 19794600, 19796400, 19798200, 19800000, 
    19801800, 19803600, 19805400, 19807200, 19809000, 19810800, 19812600, 
    19814400, 19816200, 19818000, 19819800, 19821600, 19823400, 19825200, 
    19827000, 19828800, 19830600, 19832400, 19834200, 19836000, 19837800, 
    19839600, 19841400, 19843200, 19845000, 19846800, 19848600, 19850400, 
    19852200, 19854000, 19855800, 19857600, 19859400, 19861200, 19863000, 
    19864800, 19866600, 19868400, 19870200, 19872000, 19873800, 19875600, 
    19877400, 19879200, 19881000, 19882800, 19884600, 19886400, 19888200, 
    19890000, 19891800, 19893600, 19895400, 19897200, 19899000, 19900800, 
    19902600, 19904400, 19906200, 19908000, 19909800, 19911600, 19913400, 
    19915200, 19917000, 19918800, 19920600, 19922400, 19924200, 19926000, 
    19927800, 19929600, 19931400, 19933200, 19935000, 19936800, 19938600, 
    19940400, 19942200, 19944000, 19945800, 19947600, 19949400, 19951200, 
    19953000, 19954800, 19956600, 19958400, 19960200, 19962000, 19963800, 
    19965600, 19967400, 19969200, 19971000, 19972800, 19974600, 19976400, 
    19978200, 19980000, 19981800, 19983600, 19985400, 19987200, 19989000, 
    19990800, 19992600, 19994400, 19996200, 19998000, 19999800, 20001600, 
    20003400, 20005200, 20007000, 20008800, 20010600, 20012400, 20014200, 
    20016000, 20017800, 20019600, 20021400, 20023200, 20025000, 20026800, 
    20028600, 20030400, 20032200, 20034000, 20035800, 20037600, 20039400, 
    20041200, 20043000, 20044800, 20046600, 20048400, 20050200, 20052000, 
    20053800, 20055600, 20057400, 20059200, 20061000, 20062800, 20064600, 
    20066400, 20068200, 20070000, 20071800, 20073600, 20075400, 20077200, 
    20079000, 20080800, 20082600, 20084400, 20086200, 20088000, 20089800, 
    20091600, 20093400, 20095200, 20097000, 20098800, 20100600, 20102400, 
    20104200, 20106000, 20107800, 20109600, 20111400, 20113200, 20115000, 
    20116800, 20118600, 20120400, 20122200, 20124000, 20125800, 20127600, 
    20129400, 20131200, 20133000, 20134800, 20136600, 20138400, 20140200, 
    20142000, 20143800, 20145600, 20147400, 20149200, 20151000, 20152800, 
    20154600, 20156400, 20158200, 20160000, 20161800, 20163600, 20165400, 
    20167200, 20169000, 20170800, 20172600, 20174400, 20176200, 20178000, 
    20179800, 20181600, 20183400, 20185200, 20187000, 20188800, 20190600, 
    20192400, 20194200, 20196000, 20197800, 20199600, 20201400, 20203200, 
    20205000, 20206800, 20208600, 20210400, 20212200, 20214000, 20215800, 
    20217600, 20219400, 20221200, 20223000, 20224800, 20226600, 20228400, 
    20230200, 20232000, 20233800, 20235600, 20237400, 20239200, 20241000, 
    20242800, 20244600, 20246400, 20248200, 20250000, 20251800, 20253600, 
    20255400, 20257200, 20259000, 20260800, 20262600, 20264400, 20266200, 
    20268000, 20269800, 20271600, 20273400, 20275200, 20277000, 20278800, 
    20280600, 20282400, 20284200, 20286000, 20287800, 20289600, 20291400, 
    20293200, 20295000, 20296800, 20298600, 20300400, 20302200, 20304000, 
    20305800, 20307600, 20309400, 20311200, 20313000, 20314800, 20316600, 
    20318400, 20320200, 20322000, 20323800, 20325600, 20327400, 20329200, 
    20331000, 20332800, 20334600, 20336400, 20338200, 20340000, 20341800, 
    20343600, 20345400, 20347200, 20349000, 20350800, 20352600, 20354400, 
    20356200, 20358000, 20359800, 20361600, 20363400, 20365200, 20367000, 
    20368800, 20370600, 20372400, 20374200, 20376000, 20377800, 20379600, 
    20381400, 20383200, 20385000, 20386800, 20388600, 20390400, 20392200, 
    20394000, 20395800, 20397600, 20399400, 20401200, 20403000, 20404800, 
    20406600, 20408400, 20410200, 20412000, 20413800, 20415600, 20417400, 
    20419200, 20421000, 20422800, 20424600, 20426400, 20428200, 20430000, 
    20431800, 20433600, 20435400, 20437200, 20439000, 20440800, 20442600, 
    20444400, 20446200, 20448000, 20449800, 20451600, 20453400, 20455200, 
    20457000, 20458800, 20460600, 20462400, 20464200, 20466000, 20467800, 
    20469600, 20471400, 20473200, 20475000, 20476800, 20478600, 20480400, 
    20482200, 20484000, 20485800, 20487600, 20489400, 20491200, 20493000, 
    20494800, 20496600, 20498400, 20500200, 20502000, 20503800, 20505600, 
    20507400, 20509200, 20511000, 20512800, 20514600, 20516400, 20518200, 
    20520000, 20521800, 20523600, 20525400, 20527200, 20529000, 20530800, 
    20532600, 20534400, 20536200, 20538000, 20539800, 20541600, 20543400, 
    20545200, 20547000, 20548800, 20550600, 20552400, 20554200, 20556000, 
    20557800, 20559600, 20561400, 20563200, 20565000, 20566800, 20568600, 
    20570400, 20572200, 20574000, 20575800, 20577600, 20579400, 20581200, 
    20583000, 20584800, 20586600, 20588400, 20590200, 20592000, 20593800, 
    20595600, 20597400, 20599200, 20601000, 20602800, 20604600, 20606400, 
    20608200, 20610000, 20611800, 20613600, 20615400, 20617200, 20619000, 
    20620800, 20622600, 20624400, 20626200, 20628000, 20629800, 20631600, 
    20633400, 20635200, 20637000, 20638800, 20640600, 20642400, 20644200, 
    20646000, 20647800, 20649600, 20651400, 20653200, 20655000, 20656800, 
    20658600, 20660400, 20662200, 20664000, 20665800, 20667600, 20669400, 
    20671200, 20673000, 20674800, 20676600, 20678400, 20680200, 20682000, 
    20683800, 20685600, 20687400, 20689200, 20691000, 20692800, 20694600, 
    20696400, 20698200, 20700000, 20701800, 20703600, 20705400, 20707200, 
    20709000, 20710800, 20712600, 20714400, 20716200, 20718000, 20719800, 
    20721600, 20723400, 20725200, 20727000, 20728800, 20730600, 20732400, 
    20734200, 20736000, 20737800, 20739600, 20741400, 20743200, 20745000, 
    20746800, 20748600, 20750400, 20752200, 20754000, 20755800, 20757600, 
    20759400, 20761200, 20763000, 20764800, 20766600, 20768400, 20770200, 
    20772000, 20773800, 20775600, 20777400, 20779200, 20781000, 20782800, 
    20784600, 20786400, 20788200, 20790000, 20791800, 20793600, 20795400, 
    20797200, 20799000, 20800800, 20802600, 20804400, 20806200, 20808000, 
    20809800, 20811600, 20813400, 20815200, 20817000, 20818800, 20820600, 
    20822400, 20824200, 20826000, 20827800, 20829600, 20831400, 20833200, 
    20835000, 20836800, 20838600, 20840400, 20842200, 20844000, 20845800, 
    20847600, 20849400, 20851200, 20853000, 20854800, 20856600, 20858400, 
    20860200, 20862000, 20863800, 20865600, 20867400, 20869200, 20871000, 
    20872800, 20874600, 20876400, 20878200, 20880000, 20881800, 20883600, 
    20885400, 20887200, 20889000, 20890800, 20892600, 20894400, 20896200, 
    20898000, 20899800, 20901600, 20903400, 20905200, 20907000, 20908800, 
    20910600, 20912400, 20914200, 20916000, 20917800, 20919600, 20921400, 
    20923200, 20925000, 20926800, 20928600, 20930400, 20932200, 20934000, 
    20935800, 20937600, 20939400, 20941200, 20943000, 20944800, 20946600, 
    20948400, 20950200, 20952000, 20953800, 20955600, 20957400, 20959200, 
    20961000, 20962800, 20964600, 20966400, 20968200, 20970000, 20971800, 
    20973600, 20975400, 20977200, 20979000, 20980800, 20982600, 20984400, 
    20986200, 20988000, 20989800, 20991600, 20993400, 20995200, 20997000, 
    20998800, 21000600, 21002400, 21004200, 21006000, 21007800, 21009600, 
    21011400, 21013200, 21015000, 21016800, 21018600, 21020400, 21022200, 
    21024000, 21025800, 21027600, 21029400, 21031200, 21033000, 21034800, 
    21036600, 21038400, 21040200, 21042000, 21043800, 21045600, 21047400, 
    21049200, 21051000, 21052800, 21054600, 21056400, 21058200, 21060000, 
    21061800, 21063600, 21065400, 21067200, 21069000, 21070800, 21072600, 
    21074400, 21076200, 21078000, 21079800, 21081600, 21083400, 21085200, 
    21087000, 21088800, 21090600, 21092400, 21094200, 21096000, 21097800, 
    21099600, 21101400, 21103200, 21105000, 21106800, 21108600, 21110400, 
    21112200, 21114000, 21115800, 21117600, 21119400, 21121200, 21123000, 
    21124800, 21126600, 21128400, 21130200, 21132000, 21133800, 21135600, 
    21137400, 21139200, 21141000, 21142800, 21144600, 21146400, 21148200, 
    21150000, 21151800, 21153600, 21155400, 21157200, 21159000, 21160800, 
    21162600, 21164400, 21166200, 21168000, 21169800, 21171600, 21173400, 
    21175200, 21177000, 21178800, 21180600, 21182400, 21184200, 21186000, 
    21187800, 21189600, 21191400, 21193200, 21195000, 21196800, 21198600, 
    21200400, 21202200, 21204000, 21205800, 21207600, 21209400, 21211200, 
    21213000, 21214800, 21216600, 21218400, 21220200, 21222000, 21223800, 
    21225600, 21227400, 21229200, 21231000, 21232800, 21234600, 21236400, 
    21238200, 21240000, 21241800, 21243600, 21245400, 21247200, 21249000, 
    21250800, 21252600, 21254400, 21256200, 21258000, 21259800, 21261600, 
    21263400, 21265200, 21267000, 21268800, 21270600, 21272400, 21274200, 
    21276000, 21277800, 21279600, 21281400, 21283200, 21285000, 21286800, 
    21288600, 21290400, 21292200, 21294000, 21295800, 21297600, 21299400, 
    21301200, 21303000, 21304800, 21306600, 21308400, 21310200, 21312000, 
    21313800, 21315600, 21317400, 21319200, 21321000, 21322800, 21324600, 
    21326400, 21328200, 21330000, 21331800, 21333600, 21335400, 21337200, 
    21339000, 21340800, 21342600, 21344400, 21346200, 21348000, 21349800, 
    21351600, 21353400, 21355200, 21357000, 21358800, 21360600, 21362400, 
    21364200, 21366000, 21367800, 21369600, 21371400, 21373200, 21375000, 
    21376800, 21378600, 21380400, 21382200, 21384000, 21385800, 21387600, 
    21389400, 21391200, 21393000, 21394800, 21396600, 21398400, 21400200, 
    21402000, 21403800, 21405600, 21407400, 21409200, 21411000, 21412800, 
    21414600, 21416400, 21418200, 21420000, 21421800, 21423600, 21425400, 
    21427200, 21429000, 21430800, 21432600, 21434400, 21436200, 21438000, 
    21439800, 21441600, 21443400, 21445200, 21447000, 21448800, 21450600, 
    21452400, 21454200, 21456000, 21457800, 21459600, 21461400, 21463200, 
    21465000, 21466800, 21468600, 21470400, 21472200, 21474000, 21475800, 
    21477600, 21479400, 21481200, 21483000, 21484800, 21486600, 21488400, 
    21490200, 21492000, 21493800, 21495600, 21497400, 21499200, 21501000, 
    21502800, 21504600, 21506400, 21508200, 21510000, 21511800, 21513600, 
    21515400, 21517200, 21519000, 21520800, 21522600, 21524400, 21526200, 
    21528000, 21529800, 21531600, 21533400, 21535200, 21537000, 21538800, 
    21540600, 21542400, 21544200, 21546000, 21547800, 21549600, 21551400, 
    21553200, 21555000, 21556800, 21558600, 21560400, 21562200, 21564000, 
    21565800, 21567600, 21569400, 21571200, 21573000, 21574800, 21576600, 
    21578400, 21580200, 21582000, 21583800, 21585600, 21587400, 21589200, 
    21591000, 21592800, 21594600, 21596400, 21598200, 21600000, 21601800, 
    21603600, 21605400, 21607200, 21609000, 21610800, 21612600, 21614400, 
    21616200, 21618000, 21619800, 21621600, 21623400, 21625200, 21627000, 
    21628800, 21630600, 21632400, 21634200, 21636000, 21637800, 21639600, 
    21641400, 21643200, 21645000, 21646800, 21648600, 21650400, 21652200, 
    21654000, 21655800, 21657600, 21659400, 21661200, 21663000, 21664800, 
    21666600, 21668400, 21670200, 21672000, 21673800, 21675600, 21677400, 
    21679200, 21681000, 21682800, 21684600, 21686400, 21688200, 21690000, 
    21691800, 21693600, 21695400, 21697200, 21699000, 21700800, 21702600, 
    21704400, 21706200, 21708000, 21709800, 21711600, 21713400, 21715200, 
    21717000, 21718800, 21720600, 21722400, 21724200, 21726000, 21727800, 
    21729600, 21731400, 21733200, 21735000, 21736800, 21738600, 21740400, 
    21742200, 21744000, 21745800, 21747600, 21749400, 21751200, 21753000, 
    21754800, 21756600, 21758400, 21760200, 21762000, 21763800, 21765600, 
    21767400, 21769200, 21771000, 21772800, 21774600, 21776400, 21778200, 
    21780000, 21781800, 21783600, 21785400, 21787200, 21789000, 21790800, 
    21792600, 21794400, 21796200, 21798000, 21799800, 21801600, 21803400, 
    21805200, 21807000, 21808800, 21810600, 21812400, 21814200, 21816000, 
    21817800, 21819600, 21821400, 21823200, 21825000, 21826800, 21828600, 
    21830400, 21832200, 21834000, 21835800, 21837600, 21839400, 21841200, 
    21843000, 21844800, 21846600, 21848400, 21850200, 21852000, 21853800, 
    21855600, 21857400, 21859200, 21861000, 21862800, 21864600, 21866400, 
    21868200, 21870000, 21871800, 21873600, 21875400, 21877200, 21879000, 
    21880800, 21882600, 21884400, 21886200, 21888000, 21889800, 21891600, 
    21893400, 21895200, 21897000, 21898800, 21900600, 21902400, 21904200, 
    21906000, 21907800, 21909600, 21911400, 21913200, 21915000, 21916800, 
    21918600, 21920400, 21922200, 21924000, 21925800, 21927600, 21929400, 
    21931200, 21933000, 21934800, 21936600, 21938400, 21940200, 21942000, 
    21943800, 21945600, 21947400, 21949200, 21951000, 21952800, 21954600, 
    21956400, 21958200, 21960000, 21961800, 21963600, 21965400, 21967200, 
    21969000, 21970800, 21972600, 21974400, 21976200, 21978000, 21979800, 
    21981600, 21983400, 21985200, 21987000, 21988800, 21990600, 21992400, 
    21994200, 21996000, 21997800, 21999600, 22001400, 22003200, 22005000, 
    22006800, 22008600, 22010400, 22012200, 22014000, 22015800, 22017600, 
    22019400, 22021200, 22023000, 22024800, 22026600, 22028400, 22030200, 
    22032000, 22033800, 22035600, 22037400, 22039200, 22041000, 22042800, 
    22044600, 22046400, 22048200, 22050000, 22051800, 22053600, 22055400, 
    22057200, 22059000, 22060800, 22062600, 22064400, 22066200, 22068000, 
    22069800, 22071600, 22073400, 22075200, 22077000, 22078800, 22080600, 
    22082400, 22084200, 22086000, 22087800, 22089600, 22091400, 22093200, 
    22095000, 22096800, 22098600, 22100400, 22102200, 22104000, 22105800, 
    22107600, 22109400, 22111200, 22113000, 22114800, 22116600, 22118400, 
    22120200, 22122000, 22123800, 22125600, 22127400, 22129200, 22131000, 
    22132800, 22134600, 22136400, 22138200, 22140000, 22141800, 22143600, 
    22145400, 22147200, 22149000, 22150800, 22152600, 22154400, 22156200, 
    22158000, 22159800, 22161600, 22163400, 22165200, 22167000, 22168800, 
    22170600, 22172400, 22174200, 22176000, 22177800, 22179600, 22181400, 
    22183200, 22185000, 22186800, 22188600, 22190400, 22192200, 22194000, 
    22195800, 22197600, 22199400, 22201200, 22203000, 22204800, 22206600, 
    22208400, 22210200, 22212000, 22213800, 22215600, 22217400, 22219200, 
    22221000, 22222800, 22224600, 22226400, 22228200, 22230000, 22231800, 
    22233600, 22235400, 22237200, 22239000, 22240800, 22242600, 22244400, 
    22246200, 22248000, 22249800, 22251600, 22253400, 22255200, 22257000, 
    22258800, 22260600, 22262400, 22264200, 22266000, 22267800, 22269600, 
    22271400, 22273200, 22275000, 22276800, 22278600, 22280400, 22282200, 
    22284000, 22285800, 22287600, 22289400, 22291200, 22293000, 22294800, 
    22296600, 22298400, 22300200, 22302000, 22303800, 22305600, 22307400, 
    22309200, 22311000, 22312800, 22314600, 22316400, 22318200, 22320000, 
    22321800, 22323600, 22325400, 22327200, 22329000, 22330800, 22332600, 
    22334400, 22336200, 22338000, 22339800, 22341600, 22343400, 22345200, 
    22347000, 22348800, 22350600, 22352400, 22354200, 22356000, 22357800, 
    22359600, 22361400, 22363200, 22365000, 22366800, 22368600, 22370400, 
    22372200, 22374000, 22375800, 22377600, 22379400, 22381200, 22383000, 
    22384800, 22386600, 22388400, 22390200, 22392000, 22393800, 22395600, 
    22397400, 22399200, 22401000, 22402800, 22404600, 22406400, 22408200, 
    22410000, 22411800, 22413600, 22415400, 22417200, 22419000, 22420800, 
    22422600, 22424400, 22426200, 22428000, 22429800, 22431600, 22433400, 
    22435200, 22437000, 22438800, 22440600, 22442400, 22444200, 22446000, 
    22447800, 22449600, 22451400, 22453200, 22455000, 22456800, 22458600, 
    22460400, 22462200, 22464000, 22465800, 22467600, 22469400, 22471200, 
    22473000, 22474800, 22476600, 22478400, 22480200, 22482000, 22483800, 
    22485600, 22487400, 22489200, 22491000, 22492800, 22494600, 22496400, 
    22498200, 22500000, 22501800, 22503600, 22505400, 22507200, 22509000, 
    22510800, 22512600, 22514400, 22516200, 22518000, 22519800, 22521600, 
    22523400, 22525200, 22527000, 22528800, 22530600, 22532400, 22534200, 
    22536000, 22537800, 22539600, 22541400, 22543200, 22545000, 22546800, 
    22548600, 22550400, 22552200, 22554000, 22555800, 22557600, 22559400, 
    22561200, 22563000, 22564800, 22566600, 22568400, 22570200, 22572000, 
    22573800, 22575600, 22577400, 22579200, 22581000, 22582800, 22584600, 
    22586400, 22588200, 22590000, 22591800, 22593600, 22595400, 22597200, 
    22599000, 22600800, 22602600, 22604400, 22606200, 22608000, 22609800, 
    22611600, 22613400, 22615200, 22617000, 22618800, 22620600, 22622400, 
    22624200, 22626000, 22627800, 22629600, 22631400, 22633200, 22635000, 
    22636800, 22638600, 22640400, 22642200, 22644000, 22645800, 22647600, 
    22649400, 22651200, 22653000, 22654800, 22656600, 22658400, 22660200, 
    22662000, 22663800, 22665600, 22667400, 22669200, 22671000, 22672800, 
    22674600, 22676400, 22678200, 22680000, 22681800, 22683600, 22685400, 
    22687200, 22689000, 22690800, 22692600, 22694400, 22696200, 22698000, 
    22699800, 22701600, 22703400, 22705200, 22707000, 22708800, 22710600, 
    22712400, 22714200, 22716000, 22717800, 22719600, 22721400, 22723200, 
    22725000, 22726800, 22728600, 22730400, 22732200, 22734000, 22735800, 
    22737600, 22739400, 22741200, 22743000, 22744800, 22746600, 22748400, 
    22750200, 22752000, 22753800, 22755600, 22757400, 22759200, 22761000, 
    22762800, 22764600, 22766400, 22768200, 22770000, 22771800, 22773600, 
    22775400, 22777200, 22779000, 22780800, 22782600, 22784400, 22786200, 
    22788000, 22789800, 22791600, 22793400, 22795200, 22797000, 22798800, 
    22800600, 22802400, 22804200, 22806000, 22807800, 22809600, 22811400, 
    22813200, 22815000, 22816800, 22818600, 22820400, 22822200, 22824000, 
    22825800, 22827600, 22829400, 22831200, 22833000, 22834800, 22836600, 
    22838400, 22840200, 22842000, 22843800, 22845600, 22847400, 22849200, 
    22851000, 22852800, 22854600, 22856400, 22858200, 22860000, 22861800, 
    22863600, 22865400, 22867200, 22869000, 22870800, 22872600, 22874400, 
    22876200, 22878000, 22879800, 22881600, 22883400, 22885200, 22887000, 
    22888800, 22890600, 22892400, 22894200, 22896000, 22897800, 22899600, 
    22901400, 22903200, 22905000, 22906800, 22908600, 22910400, 22912200, 
    22914000, 22915800, 22917600, 22919400, 22921200, 22923000, 22924800, 
    22926600, 22928400, 22930200, 22932000, 22933800, 22935600, 22937400, 
    22939200, 22941000, 22942800, 22944600, 22946400, 22948200, 22950000, 
    22951800, 22953600, 22955400, 22957200, 22959000, 22960800, 22962600, 
    22964400, 22966200, 22968000, 22969800, 22971600, 22973400, 22975200, 
    22977000, 22978800, 22980600, 22982400, 22984200, 22986000, 22987800, 
    22989600, 22991400, 22993200, 22995000, 22996800, 22998600, 23000400, 
    23002200, 23004000, 23005800, 23007600, 23009400, 23011200, 23013000, 
    23014800, 23016600, 23018400, 23020200, 23022000, 23023800, 23025600, 
    23027400, 23029200, 23031000, 23032800, 23034600, 23036400, 23038200, 
    23040000, 23041800, 23043600, 23045400, 23047200, 23049000, 23050800, 
    23052600, 23054400, 23056200, 23058000, 23059800, 23061600, 23063400, 
    23065200, 23067000, 23068800, 23070600, 23072400, 23074200, 23076000, 
    23077800, 23079600, 23081400, 23083200, 23085000, 23086800, 23088600, 
    23090400, 23092200, 23094000, 23095800, 23097600, 23099400, 23101200, 
    23103000, 23104800, 23106600, 23108400, 23110200, 23112000, 23113800, 
    23115600, 23117400, 23119200, 23121000, 23122800, 23124600, 23126400, 
    23128200, 23130000, 23131800, 23133600, 23135400, 23137200, 23139000, 
    23140800, 23142600, 23144400, 23146200, 23148000, 23149800, 23151600, 
    23153400, 23155200, 23157000, 23158800, 23160600, 23162400, 23164200, 
    23166000, 23167800, 23169600, 23171400, 23173200, 23175000, 23176800, 
    23178600, 23180400, 23182200, 23184000, 23185800, 23187600, 23189400, 
    23191200, 23193000, 23194800, 23196600, 23198400, 23200200, 23202000, 
    23203800, 23205600, 23207400, 23209200, 23211000, 23212800, 23214600, 
    23216400, 23218200, 23220000, 23221800, 23223600, 23225400, 23227200, 
    23229000, 23230800, 23232600, 23234400, 23236200, 23238000, 23239800, 
    23241600, 23243400, 23245200, 23247000, 23248800, 23250600, 23252400, 
    23254200, 23256000, 23257800, 23259600, 23261400, 23263200, 23265000, 
    23266800, 23268600, 23270400, 23272200, 23274000, 23275800, 23277600, 
    23279400, 23281200, 23283000, 23284800, 23286600, 23288400, 23290200, 
    23292000, 23293800, 23295600, 23297400, 23299200, 23301000, 23302800, 
    23304600, 23306400, 23308200, 23310000, 23311800, 23313600, 23315400, 
    23317200, 23319000, 23320800, 23322600, 23324400, 23326200, 23328000, 
    23329800, 23331600, 23333400, 23335200, 23337000, 23338800, 23340600, 
    23342400, 23344200, 23346000, 23347800, 23349600, 23351400, 23353200, 
    23355000, 23356800, 23358600, 23360400, 23362200, 23364000, 23365800, 
    23367600, 23369400, 23371200, 23373000, 23374800, 23376600, 23378400, 
    23380200, 23382000, 23383800, 23385600, 23387400, 23389200, 23391000, 
    23392800, 23394600, 23396400, 23398200, 23400000, 23401800, 23403600, 
    23405400, 23407200, 23409000, 23410800, 23412600, 23414400, 23416200, 
    23418000, 23419800, 23421600, 23423400, 23425200, 23427000, 23428800, 
    23430600, 23432400, 23434200, 23436000, 23437800, 23439600, 23441400, 
    23443200, 23445000, 23446800, 23448600, 23450400, 23452200, 23454000, 
    23455800, 23457600, 23459400, 23461200, 23463000, 23464800, 23466600, 
    23468400, 23470200, 23472000, 23473800, 23475600, 23477400, 23479200, 
    23481000, 23482800, 23484600, 23486400, 23488200, 23490000, 23491800, 
    23493600, 23495400, 23497200, 23499000, 23500800, 23502600, 23504400, 
    23506200, 23508000, 23509800, 23511600, 23513400, 23515200, 23517000, 
    23518800, 23520600, 23522400, 23524200, 23526000, 23527800, 23529600, 
    23531400, 23533200, 23535000, 23536800, 23538600, 23540400, 23542200, 
    23544000, 23545800, 23547600, 23549400, 23551200, 23553000, 23554800, 
    23556600, 23558400, 23560200, 23562000, 23563800, 23565600, 23567400, 
    23569200, 23571000, 23572800, 23574600, 23576400, 23578200, 23580000, 
    23581800, 23583600, 23585400, 23587200, 23589000, 23590800, 23592600, 
    23594400, 23596200, 23598000, 23599800, 23601600, 23603400, 23605200, 
    23607000, 23608800, 23610600, 23612400, 23614200, 23616000, 23617800, 
    23619600, 23621400, 23623200, 23625000, 23626800, 23628600, 23630400, 
    23632200, 23634000, 23635800, 23637600, 23639400, 23641200, 23643000, 
    23644800, 23646600, 23648400, 23650200, 23652000, 23653800, 23655600, 
    23657400, 23659200, 23661000, 23662800, 23664600, 23666400, 23668200, 
    23670000, 23671800, 23673600, 23675400, 23677200, 23679000, 23680800, 
    23682600, 23684400, 23686200, 23688000, 23689800, 23691600, 23693400, 
    23695200, 23697000, 23698800, 23700600, 23702400, 23704200, 23706000, 
    23707800, 23709600, 23711400, 23713200, 23715000, 23716800, 23718600, 
    23720400, 23722200, 23724000, 23725800, 23727600, 23729400, 23731200, 
    23733000, 23734800, 23736600, 23738400, 23740200, 23742000, 23743800, 
    23745600, 23747400, 23749200, 23751000, 23752800, 23754600, 23756400, 
    23758200, 23760000, 23761800, 23763600, 23765400, 23767200, 23769000, 
    23770800, 23772600, 23774400, 23776200, 23778000, 23779800, 23781600, 
    23783400, 23785200, 23787000, 23788800, 23790600, 23792400, 23794200, 
    23796000, 23797800, 23799600, 23801400, 23803200, 23805000, 23806800, 
    23808600, 23810400, 23812200, 23814000, 23815800, 23817600, 23819400, 
    23821200, 23823000, 23824800, 23826600, 23828400, 23830200, 23832000, 
    23833800, 23835600, 23837400, 23839200, 23841000, 23842800, 23844600, 
    23846400, 23848200, 23850000, 23851800, 23853600, 23855400, 23857200, 
    23859000, 23860800, 23862600, 23864400, 23866200, 23868000, 23869800, 
    23871600, 23873400, 23875200, 23877000, 23878800, 23880600, 23882400, 
    23884200, 23886000, 23887800, 23889600, 23891400, 23893200, 23895000, 
    23896800, 23898600, 23900400, 23902200, 23904000, 23905800, 23907600, 
    23909400, 23911200, 23913000, 23914800, 23916600, 23918400, 23920200, 
    23922000, 23923800, 23925600, 23927400, 23929200, 23931000, 23932800, 
    23934600, 23936400, 23938200, 23940000, 23941800, 23943600, 23945400, 
    23947200, 23949000, 23950800, 23952600, 23954400, 23956200, 23958000, 
    23959800, 23961600, 23963400, 23965200, 23967000, 23968800, 23970600, 
    23972400, 23974200, 23976000, 23977800, 23979600, 23981400, 23983200, 
    23985000, 23986800, 23988600, 23990400, 23992200, 23994000, 23995800, 
    23997600, 23999400, 24001200, 24003000, 24004800, 24006600, 24008400, 
    24010200, 24012000, 24013800, 24015600, 24017400, 24019200, 24021000, 
    24022800, 24024600, 24026400, 24028200, 24030000, 24031800, 24033600, 
    24035400, 24037200, 24039000, 24040800, 24042600, 24044400, 24046200, 
    24048000, 24049800, 24051600, 24053400, 24055200, 24057000, 24058800, 
    24060600, 24062400, 24064200, 24066000, 24067800, 24069600, 24071400, 
    24073200, 24075000, 24076800, 24078600, 24080400, 24082200, 24084000, 
    24085800, 24087600, 24089400, 24091200, 24093000, 24094800, 24096600, 
    24098400, 24100200, 24102000, 24103800, 24105600, 24107400, 24109200, 
    24111000, 24112800, 24114600, 24116400, 24118200, 24120000, 24121800, 
    24123600, 24125400, 24127200, 24129000, 24130800, 24132600, 24134400, 
    24136200, 24138000, 24139800, 24141600, 24143400, 24145200, 24147000, 
    24148800, 24150600, 24152400, 24154200, 24156000, 24157800, 24159600, 
    24161400, 24163200, 24165000, 24166800, 24168600, 24170400, 24172200, 
    24174000, 24175800, 24177600, 24179400, 24181200, 24183000, 24184800, 
    24186600, 24188400, 24190200, 24192000, 24193800, 24195600, 24197400, 
    24199200, 24201000, 24202800, 24204600, 24206400, 24208200, 24210000, 
    24211800, 24213600, 24215400, 24217200, 24219000, 24220800, 24222600, 
    24224400, 24226200, 24228000, 24229800, 24231600, 24233400, 24235200, 
    24237000, 24238800, 24240600, 24242400, 24244200, 24246000, 24247800, 
    24249600, 24251400, 24253200, 24255000, 24256800, 24258600, 24260400, 
    24262200, 24264000, 24265800, 24267600, 24269400, 24271200, 24273000, 
    24274800, 24276600, 24278400, 24280200, 24282000, 24283800, 24285600, 
    24287400, 24289200, 24291000, 24292800, 24294600, 24296400, 24298200, 
    24300000, 24301800, 24303600, 24305400, 24307200, 24309000, 24310800, 
    24312600, 24314400, 24316200, 24318000, 24319800, 24321600, 24323400, 
    24325200, 24327000, 24328800, 24330600, 24332400, 24334200, 24336000, 
    24337800, 24339600, 24341400, 24343200, 24345000, 24346800, 24348600, 
    24350400, 24352200, 24354000, 24355800, 24357600, 24359400, 24361200, 
    24363000, 24364800, 24366600, 24368400, 24370200, 24372000, 24373800, 
    24375600, 24377400, 24379200, 24381000, 24382800, 24384600, 24386400, 
    24388200, 24390000, 24391800, 24393600, 24395400, 24397200, 24399000, 
    24400800, 24402600, 24404400, 24406200, 24408000, 24409800, 24411600, 
    24413400, 24415200, 24417000, 24418800, 24420600, 24422400, 24424200, 
    24426000, 24427800, 24429600, 24431400, 24433200, 24435000, 24436800, 
    24438600, 24440400, 24442200, 24444000, 24445800, 24447600, 24449400, 
    24451200, 24453000, 24454800, 24456600, 24458400, 24460200, 24462000, 
    24463800, 24465600, 24467400, 24469200, 24471000, 24472800, 24474600, 
    24476400, 24478200, 24480000, 24481800, 24483600, 24485400, 24487200, 
    24489000, 24490800, 24492600, 24494400, 24496200, 24498000, 24499800, 
    24501600, 24503400, 24505200, 24507000, 24508800, 24510600, 24512400, 
    24514200, 24516000, 24517800, 24519600, 24521400, 24523200, 24525000, 
    24526800, 24528600, 24530400, 24532200, 24534000, 24535800, 24537600, 
    24539400, 24541200, 24543000, 24544800, 24546600, 24548400, 24550200, 
    24552000, 24553800, 24555600, 24557400, 24559200, 24561000, 24562800, 
    24564600, 24566400, 24568200, 24570000, 24571800, 24573600, 24575400, 
    24577200, 24579000, 24580800, 24582600, 24584400, 24586200, 24588000, 
    24589800, 24591600, 24593400, 24595200, 24597000, 24598800, 24600600, 
    24602400, 24604200, 24606000, 24607800, 24609600, 24611400, 24613200, 
    24615000, 24616800, 24618600, 24620400, 24622200, 24624000, 24625800, 
    24627600, 24629400, 24631200, 24633000, 24634800, 24636600, 24638400, 
    24640200, 24642000, 24643800, 24645600, 24647400, 24649200, 24651000, 
    24652800, 24654600, 24656400, 24658200, 24660000, 24661800, 24663600, 
    24665400, 24667200, 24669000, 24670800, 24672600, 24674400, 24676200, 
    24678000, 24679800, 24681600, 24683400, 24685200, 24687000, 24688800, 
    24690600, 24692400, 24694200, 24696000, 24697800, 24699600, 24701400, 
    24703200, 24705000, 24706800, 24708600, 24710400, 24712200, 24714000, 
    24715800, 24717600, 24719400, 24721200, 24723000, 24724800, 24726600, 
    24728400, 24730200, 24732000, 24733800, 24735600, 24737400, 24739200, 
    24741000, 24742800, 24744600, 24746400, 24748200, 24750000, 24751800, 
    24753600, 24755400, 24757200, 24759000, 24760800, 24762600, 24764400, 
    24766200, 24768000, 24769800, 24771600, 24773400, 24775200, 24777000, 
    24778800, 24780600, 24782400, 24784200, 24786000, 24787800, 24789600, 
    24791400, 24793200, 24795000, 24796800, 24798600, 24800400, 24802200, 
    24804000, 24805800, 24807600, 24809400, 24811200, 24813000, 24814800, 
    24816600, 24818400, 24820200, 24822000, 24823800, 24825600, 24827400, 
    24829200, 24831000, 24832800, 24834600, 24836400, 24838200, 24840000, 
    24841800, 24843600, 24845400, 24847200, 24849000, 24850800, 24852600, 
    24854400, 24856200, 24858000, 24859800, 24861600, 24863400, 24865200, 
    24867000, 24868800, 24870600, 24872400, 24874200, 24876000, 24877800, 
    24879600, 24881400, 24883200, 24885000, 24886800, 24888600, 24890400, 
    24892200, 24894000, 24895800, 24897600, 24899400, 24901200, 24903000, 
    24904800, 24906600, 24908400, 24910200, 24912000, 24913800, 24915600, 
    24917400, 24919200, 24921000, 24922800, 24924600, 24926400, 24928200, 
    24930000, 24931800, 24933600, 24935400, 24937200, 24939000, 24940800, 
    24942600, 24944400, 24946200, 24948000, 24949800, 24951600, 24953400, 
    24955200, 24957000, 24958800, 24960600, 24962400, 24964200, 24966000, 
    24967800, 24969600, 24971400, 24973200, 24975000, 24976800, 24978600, 
    24980400, 24982200, 24984000, 24985800, 24987600, 24989400, 24991200, 
    24993000, 24994800, 24996600, 24998400, 25000200, 25002000, 25003800, 
    25005600, 25007400, 25009200, 25011000, 25012800, 25014600, 25016400, 
    25018200, 25020000, 25021800, 25023600, 25025400, 25027200, 25029000, 
    25030800, 25032600, 25034400, 25036200, 25038000, 25039800, 25041600, 
    25043400, 25045200, 25047000, 25048800, 25050600, 25052400, 25054200, 
    25056000, 25057800, 25059600, 25061400, 25063200, 25065000, 25066800, 
    25068600, 25070400, 25072200, 25074000, 25075800, 25077600, 25079400, 
    25081200, 25083000, 25084800, 25086600, 25088400, 25090200, 25092000, 
    25093800, 25095600, 25097400, 25099200, 25101000, 25102800, 25104600, 
    25106400, 25108200, 25110000, 25111800, 25113600, 25115400, 25117200, 
    25119000, 25120800, 25122600, 25124400, 25126200, 25128000, 25129800, 
    25131600, 25133400, 25135200, 25137000, 25138800, 25140600, 25142400, 
    25144200, 25146000, 25147800, 25149600, 25151400, 25153200, 25155000, 
    25156800, 25158600, 25160400, 25162200, 25164000, 25165800, 25167600, 
    25169400, 25171200, 25173000, 25174800, 25176600, 25178400, 25180200, 
    25182000, 25183800, 25185600, 25187400, 25189200, 25191000, 25192800, 
    25194600, 25196400, 25198200, 25200000, 25201800, 25203600, 25205400, 
    25207200, 25209000, 25210800, 25212600, 25214400, 25216200, 25218000, 
    25219800, 25221600, 25223400, 25225200, 25227000, 25228800, 25230600, 
    25232400, 25234200, 25236000, 25237800, 25239600, 25241400, 25243200, 
    25245000, 25246800, 25248600, 25250400, 25252200, 25254000, 25255800, 
    25257600, 25259400, 25261200, 25263000, 25264800, 25266600, 25268400, 
    25270200, 25272000, 25273800, 25275600, 25277400, 25279200, 25281000, 
    25282800, 25284600, 25286400, 25288200, 25290000, 25291800, 25293600, 
    25295400, 25297200, 25299000, 25300800, 25302600, 25304400, 25306200, 
    25308000, 25309800, 25311600, 25313400, 25315200, 25317000, 25318800, 
    25320600, 25322400, 25324200, 25326000, 25327800, 25329600, 25331400, 
    25333200, 25335000, 25336800, 25338600, 25340400, 25342200, 25344000, 
    25345800, 25347600, 25349400, 25351200, 25353000, 25354800, 25356600, 
    25358400, 25360200, 25362000, 25363800, 25365600, 25367400, 25369200, 
    25371000, 25372800, 25374600, 25376400, 25378200, 25380000, 25381800, 
    25383600, 25385400, 25387200, 25389000, 25390800, 25392600, 25394400, 
    25396200, 25398000, 25399800, 25401600, 25403400, 25405200, 25407000, 
    25408800, 25410600, 25412400, 25414200, 25416000, 25417800, 25419600, 
    25421400, 25423200, 25425000, 25426800, 25428600, 25430400, 25432200, 
    25434000, 25435800, 25437600, 25439400, 25441200, 25443000, 25444800, 
    25446600, 25448400, 25450200, 25452000, 25453800, 25455600, 25457400, 
    25459200, 25461000, 25462800, 25464600, 25466400, 25468200, 25470000, 
    25471800, 25473600, 25475400, 25477200, 25479000, 25480800, 25482600, 
    25484400, 25486200, 25488000, 25489800, 25491600, 25493400, 25495200, 
    25497000, 25498800, 25500600, 25502400, 25504200, 25506000, 25507800, 
    25509600, 25511400, 25513200, 25515000, 25516800, 25518600, 25520400, 
    25522200, 25524000, 25525800, 25527600, 25529400, 25531200, 25533000, 
    25534800, 25536600, 25538400, 25540200, 25542000, 25543800, 25545600, 
    25547400, 25549200, 25551000, 25552800, 25554600, 25556400, 25558200, 
    25560000, 25561800, 25563600, 25565400, 25567200, 25569000, 25570800, 
    25572600, 25574400, 25576200, 25578000, 25579800, 25581600, 25583400, 
    25585200, 25587000, 25588800, 25590600, 25592400, 25594200, 25596000, 
    25597800, 25599600, 25601400, 25603200, 25605000, 25606800, 25608600, 
    25610400, 25612200, 25614000, 25615800, 25617600, 25619400, 25621200, 
    25623000, 25624800, 25626600, 25628400, 25630200, 25632000, 25633800, 
    25635600, 25637400, 25639200, 25641000, 25642800, 25644600, 25646400, 
    25648200, 25650000, 25651800, 25653600, 25655400, 25657200, 25659000, 
    25660800, 25662600, 25664400, 25666200, 25668000, 25669800, 25671600, 
    25673400, 25675200, 25677000, 25678800, 25680600, 25682400, 25684200, 
    25686000, 25687800, 25689600, 25691400, 25693200, 25695000, 25696800, 
    25698600, 25700400, 25702200, 25704000, 25705800, 25707600, 25709400, 
    25711200, 25713000, 25714800, 25716600, 25718400, 25720200, 25722000, 
    25723800, 25725600, 25727400, 25729200, 25731000, 25732800, 25734600, 
    25736400, 25738200, 25740000, 25741800, 25743600, 25745400, 25747200, 
    25749000, 25750800, 25752600, 25754400, 25756200, 25758000, 25759800, 
    25761600, 25763400, 25765200, 25767000, 25768800, 25770600, 25772400, 
    25774200, 25776000, 25777800, 25779600, 25781400, 25783200, 25785000, 
    25786800, 25788600, 25790400, 25792200, 25794000, 25795800, 25797600, 
    25799400, 25801200, 25803000, 25804800, 25806600, 25808400, 25810200, 
    25812000, 25813800, 25815600, 25817400, 25819200, 25821000, 25822800, 
    25824600, 25826400, 25828200, 25830000, 25831800, 25833600, 25835400, 
    25837200, 25839000, 25840800, 25842600, 25844400, 25846200, 25848000, 
    25849800, 25851600, 25853400, 25855200, 25857000, 25858800, 25860600, 
    25862400, 25864200, 25866000, 25867800, 25869600, 25871400, 25873200, 
    25875000, 25876800, 25878600, 25880400, 25882200, 25884000, 25885800, 
    25887600, 25889400, 25891200, 25893000, 25894800, 25896600, 25898400, 
    25900200, 25902000, 25903800, 25905600, 25907400, 25909200, 25911000, 
    25912800, 25914600, 25916400, 25918200, 25920000, 25921800, 25923600, 
    25925400, 25927200, 25929000, 25930800, 25932600, 25934400, 25936200, 
    25938000, 25939800, 25941600, 25943400, 25945200, 25947000, 25948800, 
    25950600, 25952400, 25954200, 25956000, 25957800, 25959600, 25961400, 
    25963200, 25965000, 25966800, 25968600, 25970400, 25972200, 25974000, 
    25975800, 25977600, 25979400, 25981200, 25983000, 25984800, 25986600, 
    25988400, 25990200, 25992000, 25993800, 25995600, 25997400, 25999200, 
    26001000, 26002800, 26004600, 26006400, 26008200, 26010000, 26011800, 
    26013600, 26015400, 26017200, 26019000, 26020800, 26022600, 26024400, 
    26026200, 26028000, 26029800, 26031600, 26033400, 26035200, 26037000, 
    26038800, 26040600, 26042400, 26044200, 26046000, 26047800, 26049600, 
    26051400, 26053200, 26055000, 26056800, 26058600, 26060400, 26062200, 
    26064000, 26065800, 26067600, 26069400, 26071200, 26073000, 26074800, 
    26076600, 26078400, 26080200, 26082000, 26083800, 26085600, 26087400, 
    26089200, 26091000, 26092800, 26094600, 26096400, 26098200, 26100000, 
    26101800, 26103600, 26105400, 26107200, 26109000, 26110800, 26112600, 
    26114400, 26116200, 26118000, 26119800, 26121600, 26123400, 26125200, 
    26127000, 26128800, 26130600, 26132400, 26134200, 26136000, 26137800, 
    26139600, 26141400, 26143200, 26145000, 26146800, 26148600, 26150400, 
    26152200, 26154000, 26155800, 26157600, 26159400, 26161200, 26163000, 
    26164800, 26166600, 26168400, 26170200, 26172000, 26173800, 26175600, 
    26177400, 26179200, 26181000, 26182800, 26184600, 26186400, 26188200, 
    26190000, 26191800, 26193600, 26195400, 26197200, 26199000, 26200800, 
    26202600, 26204400, 26206200, 26208000, 26209800, 26211600, 26213400, 
    26215200, 26217000, 26218800, 26220600, 26222400, 26224200, 26226000, 
    26227800, 26229600, 26231400, 26233200, 26235000, 26236800, 26238600, 
    26240400, 26242200, 26244000, 26245800, 26247600, 26249400, 26251200, 
    26253000, 26254800, 26256600, 26258400, 26260200, 26262000, 26263800, 
    26265600, 26267400, 26269200, 26271000, 26272800, 26274600, 26276400, 
    26278200, 26280000, 26281800, 26283600, 26285400, 26287200, 26289000, 
    26290800, 26292600, 26294400, 26296200, 26298000, 26299800, 26301600, 
    26303400, 26305200, 26307000, 26308800, 26310600, 26312400, 26314200, 
    26316000, 26317800, 26319600, 26321400, 26323200, 26325000, 26326800, 
    26328600, 26330400, 26332200, 26334000, 26335800, 26337600, 26339400, 
    26341200, 26343000, 26344800, 26346600, 26348400, 26350200, 26352000, 
    26353800, 26355600, 26357400, 26359200, 26361000, 26362800, 26364600, 
    26366400, 26368200, 26370000, 26371800, 26373600, 26375400, 26377200, 
    26379000, 26380800, 26382600, 26384400, 26386200, 26388000, 26389800, 
    26391600, 26393400, 26395200, 26397000, 26398800, 26400600, 26402400, 
    26404200, 26406000, 26407800, 26409600, 26411400, 26413200, 26415000, 
    26416800, 26418600, 26420400, 26422200, 26424000, 26425800, 26427600, 
    26429400, 26431200, 26433000, 26434800, 26436600, 26438400, 26440200, 
    26442000, 26443800, 26445600, 26447400, 26449200, 26451000, 26452800, 
    26454600, 26456400, 26458200, 26460000, 26461800, 26463600, 26465400, 
    26467200, 26469000, 26470800, 26472600, 26474400, 26476200, 26478000, 
    26479800, 26481600, 26483400, 26485200, 26487000, 26488800, 26490600, 
    26492400, 26494200, 26496000, 26497800, 26499600, 26501400, 26503200, 
    26505000, 26506800, 26508600, 26510400, 26512200, 26514000, 26515800, 
    26517600, 26519400, 26521200, 26523000, 26524800, 26526600, 26528400, 
    26530200, 26532000, 26533800, 26535600, 26537400, 26539200, 26541000, 
    26542800, 26544600, 26546400, 26548200, 26550000, 26551800, 26553600, 
    26555400, 26557200, 26559000, 26560800, 26562600, 26564400, 26566200, 
    26568000, 26569800, 26571600, 26573400, 26575200, 26577000, 26578800, 
    26580600, 26582400, 26584200, 26586000, 26587800, 26589600, 26591400, 
    26593200, 26595000, 26596800, 26598600, 26600400, 26602200, 26604000, 
    26605800, 26607600, 26609400, 26611200, 26613000, 26614800, 26616600, 
    26618400, 26620200, 26622000, 26623800, 26625600, 26627400, 26629200, 
    26631000, 26632800, 26634600, 26636400, 26638200, 26640000, 26641800, 
    26643600, 26645400, 26647200, 26649000, 26650800, 26652600, 26654400, 
    26656200, 26658000, 26659800, 26661600, 26663400, 26665200, 26667000, 
    26668800, 26670600, 26672400, 26674200, 26676000, 26677800, 26679600, 
    26681400, 26683200, 26685000, 26686800, 26688600, 26690400, 26692200, 
    26694000, 26695800, 26697600, 26699400, 26701200, 26703000, 26704800, 
    26706600, 26708400, 26710200, 26712000, 26713800, 26715600, 26717400, 
    26719200, 26721000, 26722800, 26724600, 26726400, 26728200, 26730000, 
    26731800, 26733600, 26735400, 26737200, 26739000, 26740800, 26742600, 
    26744400, 26746200, 26748000, 26749800, 26751600, 26753400, 26755200, 
    26757000, 26758800, 26760600, 26762400, 26764200, 26766000, 26767800, 
    26769600, 26771400, 26773200, 26775000, 26776800, 26778600, 26780400, 
    26782200, 26784000, 26785800, 26787600, 26789400, 26791200, 26793000, 
    26794800, 26796600, 26798400, 26800200, 26802000, 26803800, 26805600, 
    26807400, 26809200, 26811000, 26812800, 26814600, 26816400, 26818200, 
    26820000, 26821800, 26823600, 26825400, 26827200, 26829000, 26830800, 
    26832600, 26834400, 26836200, 26838000, 26839800, 26841600, 26843400, 
    26845200, 26847000, 26848800, 26850600, 26852400, 26854200, 26856000, 
    26857800, 26859600, 26861400, 26863200, 26865000, 26866800, 26868600, 
    26870400, 26872200, 26874000, 26875800, 26877600, 26879400, 26881200, 
    26883000, 26884800, 26886600, 26888400, 26890200, 26892000, 26893800, 
    26895600, 26897400, 26899200, 26901000, 26902800, 26904600, 26906400, 
    26908200, 26910000, 26911800, 26913600, 26915400, 26917200, 26919000, 
    26920800, 26922600, 26924400, 26926200, 26928000, 26929800, 26931600, 
    26933400, 26935200, 26937000, 26938800, 26940600, 26942400, 26944200, 
    26946000, 26947800, 26949600, 26951400, 26953200, 26955000, 26956800, 
    26958600, 26960400, 26962200, 26964000, 26965800, 26967600, 26969400, 
    26971200, 26973000, 26974800, 26976600, 26978400, 26980200, 26982000, 
    26983800, 26985600, 26987400, 26989200, 26991000, 26992800, 26994600, 
    26996400, 26998200, 27000000, 27001800, 27003600, 27005400, 27007200, 
    27009000, 27010800, 27012600, 27014400, 27016200, 27018000, 27019800, 
    27021600, 27023400, 27025200, 27027000, 27028800, 27030600, 27032400, 
    27034200, 27036000, 27037800, 27039600, 27041400, 27043200, 27045000, 
    27046800, 27048600, 27050400, 27052200, 27054000, 27055800, 27057600, 
    27059400, 27061200, 27063000, 27064800, 27066600, 27068400, 27070200, 
    27072000, 27073800, 27075600, 27077400, 27079200, 27081000, 27082800, 
    27084600, 27086400, 27088200, 27090000, 27091800, 27093600, 27095400, 
    27097200, 27099000, 27100800, 27102600, 27104400, 27106200, 27108000, 
    27109800, 27111600, 27113400, 27115200, 27117000, 27118800, 27120600, 
    27122400, 27124200, 27126000, 27127800, 27129600, 27131400, 27133200, 
    27135000, 27136800, 27138600, 27140400, 27142200, 27144000, 27145800, 
    27147600, 27149400, 27151200, 27153000, 27154800, 27156600, 27158400, 
    27160200, 27162000, 27163800, 27165600, 27167400, 27169200, 27171000, 
    27172800, 27174600, 27176400, 27178200, 27180000, 27181800, 27183600, 
    27185400, 27187200, 27189000, 27190800, 27192600, 27194400, 27196200, 
    27198000, 27199800, 27201600, 27203400, 27205200, 27207000, 27208800, 
    27210600, 27212400, 27214200, 27216000, 27217800, 27219600, 27221400, 
    27223200, 27225000, 27226800, 27228600, 27230400, 27232200, 27234000, 
    27235800, 27237600, 27239400, 27241200, 27243000, 27244800, 27246600, 
    27248400, 27250200, 27252000, 27253800, 27255600, 27257400, 27259200, 
    27261000, 27262800, 27264600, 27266400, 27268200, 27270000, 27271800, 
    27273600, 27275400, 27277200, 27279000, 27280800, 27282600, 27284400, 
    27286200, 27288000, 27289800, 27291600, 27293400, 27295200, 27297000, 
    27298800, 27300600, 27302400, 27304200, 27306000, 27307800, 27309600, 
    27311400, 27313200, 27315000, 27316800, 27318600, 27320400, 27322200, 
    27324000, 27325800, 27327600, 27329400, 27331200, 27333000, 27334800, 
    27336600, 27338400, 27340200, 27342000, 27343800, 27345600, 27347400, 
    27349200, 27351000, 27352800, 27354600, 27356400, 27358200, 27360000, 
    27361800, 27363600, 27365400, 27367200, 27369000, 27370800, 27372600, 
    27374400, 27376200, 27378000, 27379800, 27381600, 27383400, 27385200, 
    27387000, 27388800, 27390600, 27392400, 27394200, 27396000, 27397800, 
    27399600, 27401400, 27403200, 27405000, 27406800, 27408600, 27410400, 
    27412200, 27414000, 27415800, 27417600, 27419400, 27421200, 27423000, 
    27424800, 27426600, 27428400, 27430200, 27432000, 27433800, 27435600, 
    27437400, 27439200, 27441000, 27442800, 27444600, 27446400, 27448200, 
    27450000, 27451800, 27453600, 27455400, 27457200, 27459000, 27460800, 
    27462600, 27464400, 27466200, 27468000, 27469800, 27471600, 27473400, 
    27475200, 27477000, 27478800, 27480600, 27482400, 27484200, 27486000, 
    27487800, 27489600, 27491400, 27493200, 27495000, 27496800, 27498600, 
    27500400, 27502200, 27504000, 27505800, 27507600, 27509400, 27511200, 
    27513000, 27514800, 27516600, 27518400, 27520200, 27522000, 27523800, 
    27525600, 27527400, 27529200, 27531000, 27532800, 27534600, 27536400, 
    27538200, 27540000, 27541800, 27543600, 27545400, 27547200, 27549000, 
    27550800, 27552600, 27554400, 27556200, 27558000, 27559800, 27561600, 
    27563400, 27565200, 27567000, 27568800, 27570600, 27572400, 27574200, 
    27576000, 27577800, 27579600, 27581400, 27583200, 27585000, 27586800, 
    27588600, 27590400, 27592200, 27594000, 27595800, 27597600, 27599400, 
    27601200, 27603000, 27604800, 27606600, 27608400, 27610200, 27612000, 
    27613800, 27615600, 27617400, 27619200, 27621000, 27622800, 27624600, 
    27626400, 27628200, 27630000, 27631800, 27633600, 27635400, 27637200, 
    27639000, 27640800, 27642600, 27644400, 27646200, 27648000, 27649800, 
    27651600, 27653400, 27655200, 27657000, 27658800, 27660600, 27662400, 
    27664200, 27666000, 27667800, 27669600, 27671400, 27673200, 27675000, 
    27676800, 27678600, 27680400, 27682200, 27684000, 27685800, 27687600, 
    27689400, 27691200, 27693000, 27694800, 27696600, 27698400, 27700200, 
    27702000, 27703800, 27705600, 27707400, 27709200, 27711000, 27712800, 
    27714600, 27716400, 27718200, 27720000, 27721800, 27723600, 27725400, 
    27727200, 27729000, 27730800, 27732600, 27734400, 27736200, 27738000, 
    27739800, 27741600, 27743400, 27745200, 27747000, 27748800, 27750600, 
    27752400, 27754200, 27756000, 27757800, 27759600, 27761400, 27763200, 
    27765000, 27766800, 27768600, 27770400, 27772200, 27774000, 27775800, 
    27777600, 27779400, 27781200, 27783000, 27784800, 27786600, 27788400, 
    27790200, 27792000, 27793800, 27795600, 27797400, 27799200, 27801000, 
    27802800, 27804600, 27806400, 27808200, 27810000, 27811800, 27813600, 
    27815400, 27817200, 27819000, 27820800, 27822600, 27824400, 27826200, 
    27828000, 27829800, 27831600, 27833400, 27835200, 27837000, 27838800, 
    27840600, 27842400, 27844200, 27846000, 27847800, 27849600, 27851400, 
    27853200, 27855000, 27856800, 27858600, 27860400, 27862200, 27864000, 
    27865800, 27867600, 27869400, 27871200, 27873000, 27874800, 27876600, 
    27878400, 27880200, 27882000, 27883800, 27885600, 27887400, 27889200, 
    27891000, 27892800, 27894600, 27896400, 27898200, 27900000, 27901800, 
    27903600, 27905400, 27907200, 27909000, 27910800, 27912600, 27914400, 
    27916200, 27918000, 27919800, 27921600, 27923400, 27925200, 27927000, 
    27928800, 27930600, 27932400, 27934200, 27936000, 27937800, 27939600, 
    27941400, 27943200, 27945000, 27946800, 27948600, 27950400, 27952200, 
    27954000, 27955800, 27957600, 27959400, 27961200, 27963000, 27964800, 
    27966600, 27968400, 27970200, 27972000, 27973800, 27975600, 27977400, 
    27979200, 27981000, 27982800, 27984600, 27986400, 27988200, 27990000, 
    27991800, 27993600, 27995400, 27997200, 27999000, 28000800, 28002600, 
    28004400, 28006200, 28008000, 28009800, 28011600, 28013400, 28015200, 
    28017000, 28018800, 28020600, 28022400, 28024200, 28026000, 28027800, 
    28029600, 28031400, 28033200, 28035000, 28036800, 28038600, 28040400, 
    28042200, 28044000, 28045800, 28047600, 28049400, 28051200, 28053000, 
    28054800, 28056600, 28058400, 28060200, 28062000, 28063800, 28065600, 
    28067400, 28069200, 28071000, 28072800, 28074600, 28076400, 28078200, 
    28080000, 28081800, 28083600, 28085400, 28087200, 28089000, 28090800, 
    28092600, 28094400, 28096200, 28098000, 28099800, 28101600, 28103400, 
    28105200, 28107000, 28108800, 28110600, 28112400, 28114200, 28116000, 
    28117800, 28119600, 28121400, 28123200, 28125000, 28126800, 28128600, 
    28130400, 28132200, 28134000, 28135800, 28137600, 28139400, 28141200, 
    28143000, 28144800, 28146600, 28148400, 28150200, 28152000, 28153800, 
    28155600, 28157400, 28159200, 28161000, 28162800, 28164600, 28166400, 
    28168200, 28170000, 28171800, 28173600, 28175400, 28177200, 28179000, 
    28180800, 28182600, 28184400, 28186200, 28188000, 28189800, 28191600, 
    28193400, 28195200, 28197000, 28198800, 28200600, 28202400, 28204200, 
    28206000, 28207800, 28209600, 28211400, 28213200, 28215000, 28216800, 
    28218600, 28220400, 28222200, 28224000, 28225800, 28227600, 28229400, 
    28231200, 28233000, 28234800, 28236600, 28238400, 28240200, 28242000, 
    28243800, 28245600, 28247400, 28249200, 28251000, 28252800, 28254600, 
    28256400, 28258200, 28260000, 28261800, 28263600, 28265400, 28267200, 
    28269000, 28270800, 28272600, 28274400, 28276200, 28278000, 28279800, 
    28281600, 28283400, 28285200, 28287000, 28288800, 28290600, 28292400, 
    28294200, 28296000, 28297800, 28299600, 28301400, 28303200, 28305000, 
    28306800, 28308600, 28310400, 28312200, 28314000, 28315800, 28317600, 
    28319400, 28321200, 28323000, 28324800, 28326600, 28328400, 28330200, 
    28332000, 28333800, 28335600, 28337400, 28339200, 28341000, 28342800, 
    28344600, 28346400, 28348200, 28350000, 28351800, 28353600, 28355400, 
    28357200, 28359000, 28360800, 28362600, 28364400, 28366200, 28368000, 
    28369800, 28371600, 28373400, 28375200, 28377000, 28378800, 28380600, 
    28382400, 28384200, 28386000, 28387800, 28389600, 28391400, 28393200, 
    28395000, 28396800, 28398600, 28400400, 28402200, 28404000, 28405800, 
    28407600, 28409400, 28411200, 28413000, 28414800, 28416600, 28418400, 
    28420200, 28422000, 28423800, 28425600, 28427400, 28429200, 28431000, 
    28432800, 28434600, 28436400, 28438200, 28440000, 28441800, 28443600, 
    28445400, 28447200, 28449000, 28450800, 28452600, 28454400, 28456200, 
    28458000, 28459800, 28461600, 28463400, 28465200, 28467000, 28468800, 
    28470600, 28472400, 28474200, 28476000, 28477800, 28479600, 28481400, 
    28483200, 28485000, 28486800, 28488600, 28490400, 28492200, 28494000, 
    28495800, 28497600, 28499400, 28501200, 28503000, 28504800, 28506600, 
    28508400, 28510200, 28512000, 28513800, 28515600, 28517400, 28519200, 
    28521000, 28522800, 28524600, 28526400, 28528200, 28530000, 28531800, 
    28533600, 28535400, 28537200, 28539000, 28540800, 28542600, 28544400, 
    28546200, 28548000, 28549800, 28551600, 28553400, 28555200, 28557000, 
    28558800, 28560600, 28562400, 28564200, 28566000, 28567800, 28569600, 
    28571400, 28573200, 28575000, 28576800, 28578600, 28580400, 28582200, 
    28584000, 28585800, 28587600, 28589400, 28591200, 28593000, 28594800, 
    28596600, 28598400, 28600200, 28602000, 28603800, 28605600, 28607400, 
    28609200, 28611000, 28612800, 28614600, 28616400, 28618200, 28620000, 
    28621800, 28623600, 28625400, 28627200, 28629000, 28630800, 28632600, 
    28634400, 28636200, 28638000, 28639800, 28641600, 28643400, 28645200, 
    28647000, 28648800, 28650600, 28652400, 28654200, 28656000, 28657800, 
    28659600, 28661400, 28663200, 28665000, 28666800, 28668600, 28670400, 
    28672200, 28674000, 28675800, 28677600, 28679400, 28681200, 28683000, 
    28684800, 28686600, 28688400, 28690200, 28692000, 28693800, 28695600, 
    28697400, 28699200, 28701000, 28702800, 28704600, 28706400, 28708200, 
    28710000, 28711800, 28713600, 28715400, 28717200, 28719000, 28720800, 
    28722600, 28724400, 28726200, 28728000, 28729800, 28731600, 28733400, 
    28735200, 28737000, 28738800, 28740600, 28742400, 28744200, 28746000, 
    28747800, 28749600, 28751400, 28753200, 28755000, 28756800, 28758600, 
    28760400, 28762200, 28764000, 28765800, 28767600, 28769400, 28771200, 
    28773000, 28774800, 28776600, 28778400, 28780200, 28782000, 28783800, 
    28785600, 28787400, 28789200, 28791000, 28792800, 28794600, 28796400, 
    28798200, 28800000, 28801800, 28803600, 28805400, 28807200, 28809000, 
    28810800, 28812600, 28814400, 28816200, 28818000, 28819800, 28821600, 
    28823400, 28825200, 28827000, 28828800, 28830600, 28832400, 28834200, 
    28836000, 28837800, 28839600, 28841400, 28843200, 28845000, 28846800, 
    28848600, 28850400, 28852200, 28854000, 28855800, 28857600, 28859400, 
    28861200, 28863000, 28864800, 28866600, 28868400, 28870200, 28872000, 
    28873800, 28875600, 28877400, 28879200, 28881000, 28882800, 28884600, 
    28886400, 28888200, 28890000, 28891800, 28893600, 28895400, 28897200, 
    28899000, 28900800, 28902600, 28904400, 28906200, 28908000, 28909800, 
    28911600, 28913400, 28915200, 28917000, 28918800, 28920600, 28922400, 
    28924200, 28926000, 28927800, 28929600, 28931400, 28933200, 28935000, 
    28936800, 28938600, 28940400, 28942200, 28944000, 28945800, 28947600, 
    28949400, 28951200, 28953000, 28954800, 28956600, 28958400, 28960200, 
    28962000, 28963800, 28965600, 28967400, 28969200, 28971000, 28972800, 
    28974600, 28976400, 28978200, 28980000, 28981800, 28983600, 28985400, 
    28987200, 28989000, 28990800, 28992600, 28994400, 28996200, 28998000, 
    28999800, 29001600, 29003400, 29005200, 29007000, 29008800, 29010600, 
    29012400, 29014200, 29016000, 29017800, 29019600, 29021400, 29023200, 
    29025000, 29026800, 29028600, 29030400, 29032200, 29034000, 29035800, 
    29037600, 29039400, 29041200, 29043000, 29044800, 29046600, 29048400, 
    29050200, 29052000, 29053800, 29055600, 29057400, 29059200, 29061000, 
    29062800, 29064600, 29066400, 29068200, 29070000, 29071800, 29073600, 
    29075400, 29077200, 29079000, 29080800, 29082600, 29084400, 29086200, 
    29088000, 29089800, 29091600, 29093400, 29095200, 29097000, 29098800, 
    29100600, 29102400, 29104200, 29106000, 29107800, 29109600, 29111400, 
    29113200, 29115000, 29116800, 29118600, 29120400, 29122200, 29124000, 
    29125800, 29127600, 29129400, 29131200, 29133000, 29134800, 29136600, 
    29138400, 29140200, 29142000, 29143800, 29145600, 29147400, 29149200, 
    29151000, 29152800, 29154600, 29156400, 29158200, 29160000, 29161800, 
    29163600, 29165400, 29167200, 29169000, 29170800, 29172600, 29174400, 
    29176200, 29178000, 29179800, 29181600, 29183400, 29185200, 29187000, 
    29188800, 29190600, 29192400, 29194200, 29196000, 29197800, 29199600, 
    29201400, 29203200, 29205000, 29206800, 29208600, 29210400, 29212200, 
    29214000, 29215800, 29217600, 29219400, 29221200, 29223000, 29224800, 
    29226600, 29228400, 29230200, 29232000, 29233800, 29235600, 29237400, 
    29239200, 29241000, 29242800, 29244600, 29246400, 29248200, 29250000, 
    29251800, 29253600, 29255400, 29257200, 29259000, 29260800, 29262600, 
    29264400, 29266200, 29268000, 29269800, 29271600, 29273400, 29275200, 
    29277000, 29278800, 29280600, 29282400, 29284200, 29286000, 29287800, 
    29289600, 29291400, 29293200, 29295000, 29296800, 29298600, 29300400, 
    29302200, 29304000, 29305800, 29307600, 29309400, 29311200, 29313000, 
    29314800, 29316600, 29318400, 29320200, 29322000, 29323800, 29325600, 
    29327400, 29329200, 29331000, 29332800, 29334600, 29336400, 29338200, 
    29340000, 29341800, 29343600, 29345400, 29347200, 29349000, 29350800, 
    29352600, 29354400, 29356200, 29358000, 29359800, 29361600, 29363400, 
    29365200, 29367000, 29368800, 29370600, 29372400, 29374200, 29376000, 
    29377800, 29379600, 29381400, 29383200, 29385000, 29386800, 29388600, 
    29390400, 29392200, 29394000, 29395800, 29397600, 29399400, 29401200, 
    29403000, 29404800, 29406600, 29408400, 29410200, 29412000, 29413800, 
    29415600, 29417400, 29419200, 29421000, 29422800, 29424600, 29426400, 
    29428200, 29430000, 29431800, 29433600, 29435400, 29437200, 29439000, 
    29440800, 29442600, 29444400, 29446200, 29448000, 29449800, 29451600, 
    29453400, 29455200, 29457000, 29458800, 29460600, 29462400, 29464200, 
    29466000, 29467800, 29469600, 29471400, 29473200, 29475000, 29476800, 
    29478600, 29480400, 29482200, 29484000, 29485800, 29487600, 29489400, 
    29491200, 29493000, 29494800, 29496600, 29498400, 29500200, 29502000, 
    29503800, 29505600, 29507400, 29509200, 29511000, 29512800, 29514600, 
    29516400, 29518200, 29520000, 29521800, 29523600, 29525400, 29527200, 
    29529000, 29530800, 29532600, 29534400, 29536200, 29538000, 29539800, 
    29541600, 29543400, 29545200, 29547000, 29548800, 29550600, 29552400, 
    29554200, 29556000, 29557800, 29559600, 29561400, 29563200, 29565000, 
    29566800, 29568600, 29570400, 29572200, 29574000, 29575800, 29577600, 
    29579400, 29581200, 29583000, 29584800, 29586600, 29588400, 29590200, 
    29592000, 29593800, 29595600, 29597400, 29599200, 29601000, 29602800, 
    29604600, 29606400, 29608200, 29610000, 29611800, 29613600, 29615400, 
    29617200, 29619000, 29620800, 29622600, 29624400, 29626200, 29628000, 
    29629800, 29631600, 29633400, 29635200, 29637000, 29638800, 29640600, 
    29642400, 29644200, 29646000, 29647800, 29649600, 29651400, 29653200, 
    29655000, 29656800, 29658600, 29660400, 29662200, 29664000, 29665800, 
    29667600, 29669400, 29671200, 29673000, 29674800, 29676600, 29678400, 
    29680200, 29682000, 29683800, 29685600, 29687400, 29689200, 29691000, 
    29692800, 29694600, 29696400, 29698200, 29700000, 29701800, 29703600, 
    29705400, 29707200, 29709000, 29710800, 29712600, 29714400, 29716200, 
    29718000, 29719800, 29721600, 29723400, 29725200, 29727000, 29728800, 
    29730600, 29732400, 29734200, 29736000, 29737800, 29739600, 29741400, 
    29743200, 29745000, 29746800, 29748600, 29750400, 29752200, 29754000, 
    29755800, 29757600, 29759400, 29761200, 29763000, 29764800, 29766600, 
    29768400, 29770200, 29772000, 29773800, 29775600, 29777400, 29779200, 
    29781000, 29782800, 29784600, 29786400, 29788200, 29790000, 29791800, 
    29793600, 29795400, 29797200, 29799000, 29800800, 29802600, 29804400, 
    29806200, 29808000, 29809800, 29811600, 29813400, 29815200, 29817000, 
    29818800, 29820600, 29822400, 29824200, 29826000, 29827800, 29829600, 
    29831400, 29833200, 29835000, 29836800, 29838600, 29840400, 29842200, 
    29844000, 29845800, 29847600, 29849400, 29851200, 29853000, 29854800, 
    29856600, 29858400, 29860200, 29862000, 29863800, 29865600, 29867400, 
    29869200, 29871000, 29872800, 29874600, 29876400, 29878200, 29880000, 
    29881800, 29883600, 29885400, 29887200, 29889000, 29890800, 29892600, 
    29894400, 29896200, 29898000, 29899800, 29901600, 29903400, 29905200, 
    29907000, 29908800, 29910600, 29912400, 29914200, 29916000, 29917800, 
    29919600, 29921400, 29923200, 29925000, 29926800, 29928600, 29930400, 
    29932200, 29934000, 29935800, 29937600, 29939400, 29941200, 29943000, 
    29944800, 29946600, 29948400, 29950200, 29952000, 29953800, 29955600, 
    29957400, 29959200, 29961000, 29962800, 29964600, 29966400, 29968200, 
    29970000, 29971800, 29973600, 29975400, 29977200, 29979000, 29980800, 
    29982600, 29984400, 29986200, 29988000, 29989800, 29991600, 29993400, 
    29995200, 29997000, 29998800, 30000600, 30002400, 30004200, 30006000, 
    30007800, 30009600, 30011400, 30013200, 30015000, 30016800, 30018600, 
    30020400, 30022200, 30024000, 30025800, 30027600, 30029400, 30031200, 
    30033000, 30034800, 30036600, 30038400, 30040200, 30042000, 30043800, 
    30045600, 30047400, 30049200, 30051000, 30052800, 30054600, 30056400, 
    30058200, 30060000, 30061800, 30063600, 30065400, 30067200, 30069000, 
    30070800, 30072600, 30074400, 30076200, 30078000, 30079800, 30081600, 
    30083400, 30085200, 30087000, 30088800, 30090600, 30092400, 30094200, 
    30096000, 30097800, 30099600, 30101400, 30103200, 30105000, 30106800, 
    30108600, 30110400, 30112200, 30114000, 30115800, 30117600, 30119400, 
    30121200, 30123000, 30124800, 30126600, 30128400, 30130200, 30132000, 
    30133800, 30135600, 30137400, 30139200, 30141000, 30142800, 30144600, 
    30146400, 30148200, 30150000, 30151800, 30153600, 30155400, 30157200, 
    30159000, 30160800, 30162600, 30164400, 30166200, 30168000, 30169800, 
    30171600, 30173400, 30175200, 30177000, 30178800, 30180600, 30182400, 
    30184200, 30186000, 30187800, 30189600, 30191400, 30193200, 30195000, 
    30196800, 30198600, 30200400, 30202200, 30204000, 30205800, 30207600, 
    30209400, 30211200, 30213000, 30214800, 30216600, 30218400, 30220200, 
    30222000, 30223800, 30225600, 30227400, 30229200, 30231000, 30232800, 
    30234600, 30236400, 30238200, 30240000, 30241800, 30243600, 30245400, 
    30247200, 30249000, 30250800, 30252600, 30254400, 30256200, 30258000, 
    30259800, 30261600, 30263400, 30265200, 30267000, 30268800, 30270600, 
    30272400, 30274200, 30276000, 30277800, 30279600, 30281400, 30283200, 
    30285000, 30286800, 30288600, 30290400, 30292200, 30294000, 30295800, 
    30297600, 30299400, 30301200, 30303000, 30304800, 30306600, 30308400, 
    30310200, 30312000, 30313800, 30315600, 30317400, 30319200, 30321000, 
    30322800, 30324600, 30326400, 30328200, 30330000, 30331800, 30333600, 
    30335400, 30337200, 30339000, 30340800, 30342600, 30344400, 30346200, 
    30348000, 30349800, 30351600, 30353400, 30355200, 30357000, 30358800, 
    30360600, 30362400, 30364200, 30366000, 30367800, 30369600, 30371400, 
    30373200, 30375000, 30376800, 30378600, 30380400, 30382200, 30384000, 
    30385800, 30387600, 30389400, 30391200, 30393000, 30394800, 30396600, 
    30398400, 30400200, 30402000, 30403800, 30405600, 30407400, 30409200, 
    30411000, 30412800, 30414600, 30416400, 30418200, 30420000, 30421800, 
    30423600, 30425400, 30427200, 30429000, 30430800, 30432600, 30434400, 
    30436200, 30438000, 30439800, 30441600, 30443400, 30445200, 30447000, 
    30448800, 30450600, 30452400, 30454200, 30456000, 30457800, 30459600, 
    30461400, 30463200, 30465000, 30466800, 30468600, 30470400, 30472200, 
    30474000, 30475800, 30477600, 30479400, 30481200, 30483000, 30484800, 
    30486600, 30488400, 30490200, 30492000, 30493800, 30495600, 30497400, 
    30499200, 30501000, 30502800, 30504600, 30506400, 30508200, 30510000, 
    30511800, 30513600, 30515400, 30517200, 30519000, 30520800, 30522600, 
    30524400, 30526200, 30528000, 30529800, 30531600, 30533400, 30535200, 
    30537000, 30538800, 30540600, 30542400, 30544200, 30546000, 30547800, 
    30549600, 30551400, 30553200, 30555000, 30556800, 30558600, 30560400, 
    30562200, 30564000, 30565800, 30567600, 30569400, 30571200, 30573000, 
    30574800, 30576600, 30578400, 30580200, 30582000, 30583800, 30585600, 
    30587400, 30589200, 30591000, 30592800, 30594600, 30596400, 30598200, 
    30600000, 30601800, 30603600, 30605400, 30607200, 30609000, 30610800, 
    30612600, 30614400, 30616200, 30618000, 30619800, 30621600, 30623400, 
    30625200, 30627000, 30628800, 30630600, 30632400, 30634200, 30636000, 
    30637800, 30639600, 30641400, 30643200, 30645000, 30646800, 30648600, 
    30650400, 30652200, 30654000, 30655800, 30657600, 30659400, 30661200, 
    30663000, 30664800, 30666600, 30668400, 30670200, 30672000, 30673800, 
    30675600, 30677400, 30679200, 30681000, 30682800, 30684600, 30686400, 
    30688200, 30690000, 30691800, 30693600, 30695400, 30697200, 30699000, 
    30700800, 30702600, 30704400, 30706200, 30708000, 30709800, 30711600, 
    30713400, 30715200, 30717000, 30718800, 30720600, 30722400, 30724200, 
    30726000, 30727800, 30729600, 30731400, 30733200, 30735000, 30736800, 
    30738600, 30740400, 30742200, 30744000, 30745800, 30747600, 30749400, 
    30751200, 30753000, 30754800, 30756600, 30758400, 30760200, 30762000, 
    30763800, 30765600, 30767400, 30769200, 30771000, 30772800, 30774600, 
    30776400, 30778200, 30780000, 30781800, 30783600, 30785400, 30787200, 
    30789000, 30790800, 30792600, 30794400, 30796200, 30798000, 30799800, 
    30801600, 30803400, 30805200, 30807000, 30808800, 30810600, 30812400, 
    30814200, 30816000, 30817800, 30819600, 30821400, 30823200, 30825000, 
    30826800, 30828600, 30830400, 30832200, 30834000, 30835800, 30837600, 
    30839400, 30841200, 30843000, 30844800, 30846600, 30848400, 30850200, 
    30852000, 30853800, 30855600, 30857400, 30859200, 30861000, 30862800, 
    30864600, 30866400, 30868200, 30870000, 30871800, 30873600, 30875400, 
    30877200, 30879000, 30880800, 30882600, 30884400, 30886200, 30888000, 
    30889800, 30891600, 30893400, 30895200, 30897000, 30898800, 30900600, 
    30902400, 30904200, 30906000, 30907800, 30909600, 30911400, 30913200, 
    30915000, 30916800, 30918600, 30920400, 30922200, 30924000, 30925800, 
    30927600, 30929400, 30931200, 30933000, 30934800, 30936600, 30938400, 
    30940200, 30942000, 30943800, 30945600, 30947400, 30949200, 30951000, 
    30952800, 30954600, 30956400, 30958200, 30960000, 30961800, 30963600, 
    30965400, 30967200, 30969000, 30970800, 30972600, 30974400, 30976200, 
    30978000, 30979800, 30981600, 30983400, 30985200, 30987000, 30988800, 
    30990600, 30992400, 30994200, 30996000, 30997800, 30999600, 31001400, 
    31003200, 31005000, 31006800, 31008600, 31010400, 31012200, 31014000, 
    31015800, 31017600, 31019400, 31021200, 31023000, 31024800, 31026600, 
    31028400, 31030200, 31032000, 31033800, 31035600, 31037400, 31039200, 
    31041000, 31042800, 31044600, 31046400, 31048200, 31050000, 31051800, 
    31053600, 31055400, 31057200, 31059000, 31060800, 31062600, 31064400, 
    31066200, 31068000, 31069800, 31071600, 31073400, 31075200, 31077000, 
    31078800, 31080600, 31082400, 31084200, 31086000, 31087800, 31089600, 
    31091400, 31093200, 31095000, 31096800, 31098600, 31100400, 31102200, 
    31104000, 31105800, 31107600, 31109400, 31111200, 31113000, 31114800, 
    31116600, 31118400, 31120200, 31122000, 31123800, 31125600, 31127400, 
    31129200, 31131000, 31132800, 31134600, 31136400, 31138200, 31140000, 
    31141800, 31143600, 31145400, 31147200, 31149000, 31150800, 31152600, 
    31154400, 31156200, 31158000, 31159800, 31161600, 31163400, 31165200, 
    31167000, 31168800, 31170600, 31172400, 31174200, 31176000, 31177800, 
    31179600, 31181400, 31183200, 31185000, 31186800, 31188600, 31190400, 
    31192200, 31194000, 31195800, 31197600, 31199400, 31201200, 31203000, 
    31204800, 31206600, 31208400, 31210200, 31212000, 31213800, 31215600, 
    31217400, 31219200, 31221000, 31222800, 31224600, 31226400, 31228200, 
    31230000, 31231800, 31233600, 31235400, 31237200, 31239000, 31240800, 
    31242600, 31244400, 31246200, 31248000, 31249800, 31251600, 31253400, 
    31255200, 31257000, 31258800, 31260600, 31262400, 31264200, 31266000, 
    31267800, 31269600, 31271400, 31273200, 31275000, 31276800, 31278600, 
    31280400, 31282200, 31284000, 31285800, 31287600, 31289400, 31291200, 
    31293000, 31294800, 31296600, 31298400, 31300200, 31302000, 31303800, 
    31305600, 31307400, 31309200, 31311000, 31312800, 31314600, 31316400, 
    31318200, 31320000, 31321800, 31323600, 31325400, 31327200, 31329000, 
    31330800, 31332600, 31334400, 31336200, 31338000, 31339800, 31341600, 
    31343400, 31345200, 31347000, 31348800, 31350600, 31352400, 31354200, 
    31356000, 31357800, 31359600, 31361400, 31363200, 31365000, 31366800, 
    31368600, 31370400, 31372200, 31374000, 31375800, 31377600, 31379400, 
    31381200, 31383000, 31384800, 31386600, 31388400, 31390200, 31392000, 
    31393800, 31395600, 31397400, 31399200, 31401000, 31402800, 31404600, 
    31406400, 31408200, 31410000, 31411800, 31413600, 31415400, 31417200, 
    31419000, 31420800, 31422600, 31424400, 31426200, 31428000, 31429800, 
    31431600, 31433400, 31435200, 31437000, 31438800, 31440600, 31442400, 
    31444200, 31446000, 31447800, 31449600, 31451400, 31453200, 31455000, 
    31456800, 31458600, 31460400, 31462200, 31464000, 31465800, 31467600, 
    31469400, 31471200, 31473000, 31474800, 31476600, 31478400, 31480200, 
    31482000, 31483800, 31485600, 31487400, 31489200, 31491000, 31492800, 
    31494600, 31496400, 31498200, 31500000, 31501800, 31503600, 31505400, 
    31507200, 31509000, 31510800, 31512600, 31514400, 31516200, 31518000, 
    31519800, 31521600, 31523400, 31525200, 31527000, 31528800, 31530600, 
    31532400, 31534200 ;

 z = 4 ;

 y = 1 ;

 x = 1 ;

 latitude =
  52.16658 ;

 longitude =
  5.74356 ;

 SWdown =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.3,
  36.5,
  89.5,
  142.3,
  191.4,
  227.9,
  255.3,
  269.5,
  270.9,
  257.7,
  233.1,
  195.8,
  152.5,
  107.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.1,
  31.8,
  93.5,
  157.9,
  200.7,
  218.1,
  249.1,
  278.9,
  295.9,
  289.9,
  259.5,
  217.3,
  168.4,
  114.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  6.2,
  18,
  38.8,
  49.2,
  71.5,
  75,
  88.9,
  76,
  107.3,
  113.2,
  110.5,
  100.3,
  32,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  6.1,
  15.1,
  35.6,
  54,
  68.4,
  63.2,
  69.9,
  66.5,
  71.2,
  70.5,
  42.8,
  30,
  27.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.8,
  12.6,
  32.4,
  43.7,
  61.9,
  68.8,
  64.1,
  72.8,
  78.6,
  97.5,
  110,
  144.5,
  169.9,
  117.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.5,
  4.6,
  13.1,
  20,
  35.5,
  47.7,
  84.5,
  153.9,
  227.6,
  333,
  315.3,
  261.1,
  206.2,
  147.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  4.3,
  11.2,
  20.2,
  37.3,
  77.6,
  78.4,
  88.2,
  79.4,
  95.7,
  97.7,
  126.4,
  89.2,
  79,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.5,
  8,
  18,
  29.7,
  39.9,
  42.6,
  46,
  50.7,
  66,
  78,
  69.7,
  53,
  51.8,
  39.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  7.2,
  17.7,
  30.2,
  42.5,
  58.8,
  77.7,
  80.7,
  79.5,
  78.6,
  64.8,
  65.2,
  59.1,
  47,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  4.1,
  8.9,
  15.4,
  29.5,
  43.2,
  43,
  77.6,
  84.2,
  87.3,
  60.6,
  52.2,
  34.5,
  17.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.1,
  6.7,
  16.3,
  25.3,
  31.2,
  35.2,
  40.4,
  49.3,
  56.3,
  64.1,
  67,
  64.8,
  53.8,
  41.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.1,
  14.2,
  23.3,
  33.6,
  47.8,
  65.2,
  43.9,
  74,
  101.3,
  82.9,
  68.3,
  46.6,
  38.1,
  33.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.5,
  14.7,
  43.5,
  52.3,
  82.2,
  215.6,
  244.2,
  276.2,
  240,
  231.4,
  242,
  232.5,
  166.5,
  121.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.4,
  41.3,
  67.1,
  122.4,
  193.1,
  167.9,
  199.7,
  191.4,
  232.2,
  267.5,
  239.4,
  240.2,
  201.5,
  159.7,
  118.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.6,
  33.7,
  77.7,
  125.6,
  171.5,
  206.8,
  235,
  256,
  263.8,
  264.1,
  247.6,
  221,
  184.7,
  140,
  88.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.8,
  39.8,
  88.6,
  136.7,
  181.8,
  218.6,
  247.1,
  266.3,
  275.2,
  273.3,
  256.3,
  231.3,
  194.8,
  151.3,
  98.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.8,
  37.7,
  83.1,
  130.7,
  175.7,
  212.6,
  241.3,
  262.4,
  269.9,
  264.8,
  251,
  226.5,
  191.2,
  148.1,
  89.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  5.6,
  14.6,
  17.9,
  24.6,
  22.1,
  24.3,
  34.6,
  27.5,
  26.8,
  32.4,
  29.6,
  22.6,
  19.2,
  11.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.4,
  7.2,
  22.1,
  37.1,
  44.7,
  38.5,
  31.3,
  21.6,
  22.6,
  24.4,
  30,
  27.8,
  52.1,
  26.6,
  42.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.7,
  5.5,
  11.1,
  24,
  37.8,
  57.5,
  87.3,
  159.4,
  175.8,
  130.8,
  134.3,
  85.2,
  53.6,
  35.5,
  35.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.5,
  20.8,
  49,
  100.2,
  99.2,
  92.7,
  79.3,
  76.3,
  79.5,
  83.7,
  61.8,
  55.5,
  47.8,
  42.1,
  20.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.5,
  18.1,
  49,
  63.3,
  121.5,
  121.3,
  128.8,
  77.8,
  110,
  135.9,
  191.4,
  143.5,
  136.4,
  62.8,
  105.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.2,
  34.4,
  58.7,
  58.3,
  41.5,
  68.7,
  98.1,
  233.8,
  120.1,
  65.3,
  82.1,
  66.1,
  69.4,
  120.3,
  102.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.2,
  17.2,
  36.8,
  82.6,
  140.2,
  149.1,
  134.2,
  178.2,
  183.9,
  212.4,
  198.3,
  198.3,
  205.4,
  167,
  112,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.4,
  10,
  24.9,
  67.8,
  133.8,
  244.4,
  256.2,
  281.3,
  298,
  305.1,
  278.2,
  240,
  214.8,
  211.1,
  192.6,
  112.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.2,
  9.5,
  15.8,
  24.5,
  29.1,
  34.8,
  41.3,
  56.6,
  55.8,
  54.6,
  38.2,
  31.7,
  26.6,
  20.4,
  16.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  10.7,
  33.6,
  42.4,
  52.4,
  73.7,
  98.4,
  119.7,
  93.6,
  97.2,
  100.2,
  79.4,
  74.5,
  56.2,
  44.3,
  31.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.6,
  4.2,
  12.3,
  35.5,
  57.3,
  69.4,
  87,
  93.7,
  98.7,
  91.8,
  83.1,
  69.3,
  47.7,
  44.4,
  45.8,
  30.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  5.4,
  16.5,
  28.3,
  38.8,
  57.1,
  58.1,
  59.3,
  91.8,
  95,
  71.8,
  77.8,
  55,
  54.3,
  47.1,
  29.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  9.7,
  12.4,
  14,
  21.3,
  31,
  39.7,
  48.5,
  48.8,
  53.4,
  49.9,
  48.4,
  41.4,
  33.8,
  27.6,
  20.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.7,
  11.8,
  20.8,
  26.4,
  46.5,
  32,
  46.5,
  62.2,
  75.3,
  67.9,
  96.1,
  106,
  119.1,
  136,
  114.4,
  106.9,
  20.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.4,
  7.4,
  19,
  33.8,
  58.6,
  75.3,
  93.5,
  112.1,
  122.3,
  121.6,
  124.8,
  138.9,
  172.3,
  160.2,
  103.2,
  70.1,
  34.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.2,
  18.6,
  43.5,
  92.4,
  199.5,
  251.6,
  297.2,
  140,
  186.6,
  260.9,
  312,
  214.2,
  153,
  197,
  98.8,
  51.3,
  18.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.4,
  12.8,
  30.5,
  48.5,
  70.3,
  87.3,
  106.6,
  115.9,
  109,
  108.1,
  101.7,
  97.8,
  107.9,
  85.2,
  54.2,
  41.8,
  34.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.7,
  12,
  20,
  25,
  30.4,
  31.2,
  33.1,
  35.9,
  35,
  25.9,
  35.4,
  31.8,
  22.7,
  18.3,
  18.8,
  12.3,
  7.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  8,
  32.8,
  48.8,
  218,
  230.7,
  263.2,
  267.3,
  322,
  295.3,
  235.1,
  260.9,
  184.2,
  122.7,
  110.2,
  68.9,
  33.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.2,
  6.9,
  16.8,
  30.7,
  53.1,
  75.7,
  74.7,
  80.1,
  168.2,
  172.2,
  188.6,
  244.7,
  165.1,
  174.3,
  96.8,
  52.2,
  54.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.5,
  6.7,
  21,
  65.6,
  83,
  88.6,
  117.8,
  148.6,
  187.2,
  200.8,
  283.9,
  97.5,
  73,
  51.7,
  63.8,
  31.4,
  24.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.4,
  32.4,
  72.6,
  94.1,
  136.2,
  106,
  125,
  304.5,
  269.8,
  269.2,
  265.4,
  205.3,
  261.3,
  275.6,
  212,
  126.8,
  94.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.3,
  36.3,
  74.6,
  128.2,
  173.4,
  139.7,
  89.3,
  44.5,
  58.7,
  138.3,
  137,
  277.8,
  267.6,
  191,
  100.4,
  43.4,
  25.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.9,
  14.1,
  41.4,
  77.4,
  45.1,
  99.1,
  95.3,
  104.7,
  126.3,
  95,
  39.8,
  41,
  80.1,
  28.2,
  20.1,
  12.4,
  11,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  8.1,
  49,
  105.5,
  114.1,
  164.5,
  194.4,
  204,
  319.8,
  165.2,
  92.1,
  141.9,
  154.5,
  96.1,
  96.7,
  105,
  81.7,
  58.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.3,
  7.3,
  8.4,
  17.8,
  17,
  18.8,
  23,
  18.3,
  42.8,
  34.2,
  24.4,
  26,
  24.8,
  18,
  24.5,
  24.4,
  11.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  4.8,
  7.1,
  13.7,
  30,
  115.8,
  137.3,
  208.3,
  170.7,
  172.1,
  111.6,
  85,
  64.7,
  33.7,
  50.5,
  30.7,
  15.7,
  17.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  16.7,
  61.1,
  108.9,
  183.6,
  243.6,
  271.9,
  337.1,
  383.3,
  408.7,
  461.9,
  325.9,
  409.6,
  255.3,
  189.4,
  176.2,
  92.6,
  185.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.9,
  11.1,
  29.1,
  68.4,
  140.4,
  221.4,
  263.8,
  307.7,
  326.5,
  441.8,
  345.5,
  247.6,
  239.9,
  184.9,
  138.8,
  272,
  292.8,
  192.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.5,
  37.2,
  67.8,
  85.9,
  117.3,
  177.9,
  125.6,
  172.3,
  179.3,
  163.7,
  226.6,
  223.1,
  213.3,
  247.8,
  240.5,
  153.2,
  114.9,
  76,
  46.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.9,
  11.7,
  20.2,
  30.1,
  38.3,
  38.6,
  47.2,
  54.3,
  58.7,
  52.9,
  155.3,
  161.8,
  123.9,
  217.7,
  168.9,
  128.5,
  89.6,
  30.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.4,
  5.2,
  13.1,
  16.6,
  19.4,
  151.4,
  216.6,
  87.8,
  238.3,
  107,
  280.3,
  197,
  217.3,
  180.5,
  174.8,
  144.2,
  94.2,
  59.6,
  84.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.9,
  30.9,
  82.9,
  128.7,
  178.2,
  276.2,
  317.6,
  335.8,
  279.8,
  202.3,
  174.6,
  159.9,
  108.3,
  66.9,
  65.3,
  75.1,
  68.9,
  83.2,
  40.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4,
  33.6,
  86.7,
  153,
  216,
  266.3,
  321.8,
  365.4,
  297.3,
  281.2,
  253.6,
  316.9,
  290,
  266.4,
  174.6,
  148.7,
  106.3,
  73.1,
  45.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.6,
  4.2,
  10.1,
  16.1,
  30.1,
  34.1,
  33.8,
  26.1,
  25.1,
  24.4,
  26.9,
  31.5,
  50.7,
  38.9,
  47.9,
  74.9,
  59.6,
  71.3,
  25.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.6,
  6.4,
  15.2,
  29.7,
  31.8,
  48.3,
  49.9,
  43.1,
  58.8,
  77.9,
  53.7,
  83.3,
  114.8,
  146.4,
  125.3,
  93.5,
  65.7,
  50.7,
  20.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.6,
  19.8,
  41.1,
  48.3,
  92.4,
  142.5,
  181.5,
  271.9,
  335.1,
  311.7,
  355.5,
  227.9,
  270.6,
  221.5,
  154,
  116.4,
  128.9,
  69.2,
  27,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.2,
  4.7,
  5.2,
  8.5,
  60.3,
  74.5,
  73.1,
  56.2,
  79.4,
  135.1,
  113,
  58.2,
  37,
  46.9,
  34.1,
  76.2,
  70.6,
  206,
  48.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  8.2,
  36.3,
  53.6,
  65.1,
  27.8,
  78.6,
  253.9,
  240,
  395.7,
  246.8,
  252.2,
  197.5,
  127.5,
  148.1,
  123.2,
  105,
  85.2,
  77.5,
  53.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  20.7,
  34.6,
  76.7,
  46.6,
  49.8,
  132.9,
  113.6,
  68.6,
  140.4,
  149.8,
  120.3,
  34.3,
  71,
  188.3,
  144.1,
  90.5,
  33.5,
  68.7,
  50.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  18.2,
  57.3,
  129.4,
  179.5,
  151.7,
  52.8,
  111.3,
  137.8,
  206.1,
  219.9,
  195.8,
  165.3,
  172.7,
  177.2,
  124.2,
  121,
  150.5,
  134.8,
  69.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  12.4,
  46.8,
  83.4,
  152.5,
  236.6,
  297.8,
  295,
  229.6,
  260.1,
  372.1,
  312.7,
  457.9,
  354,
  352.5,
  274.8,
  248.1,
  233.6,
  139.9,
  79.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  19.7,
  92.2,
  178.6,
  154.8,
  242.5,
  335.9,
  392.3,
  439.5,
  472.5,
  469.5,
  427,
  422.1,
  338.3,
  284.7,
  282.9,
  293.5,
  296,
  196.1,
  149.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  7.5,
  32.3,
  41.5,
  58.8,
  44.2,
  38.8,
  90.7,
  210.2,
  222.4,
  54.6,
  31,
  34.3,
  26.7,
  20.4,
  18.2,
  19.2,
  20.3,
  30.7,
  29.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  13.3,
  67.6,
  91.5,
  151.9,
  155,
  263.7,
  391.9,
  451.4,
  475.6,
  498,
  490.9,
  518.3,
  377.9,
  384,
  343.7,
  212.5,
  152.2,
  104.5,
  71.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.5,
  25.6,
  83.7,
  152.6,
  223.3,
  284.2,
  319.9,
  353.1,
  230.5,
  231.1,
  202.8,
  183,
  233.4,
  320,
  237.1,
  259.4,
  168.8,
  219.6,
  160.7,
  84.6,
  46.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.8,
  9.2,
  14,
  23.1,
  31.4,
  93.6,
  163.3,
  215.8,
  143.8,
  98.3,
  398.5,
  207.5,
  201.2,
  204,
  298.6,
  377.6,
  309.7,
  232.9,
  224.6,
  159.4,
  92.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  8.7,
  19.7,
  31.2,
  52.6,
  162.5,
  339.3,
  455.1,
  427.3,
  477.4,
  352,
  612.8,
  564.7,
  428,
  421.3,
  350.8,
  360,
  296.5,
  101.6,
  61.4,
  50.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.2,
  25,
  44.6,
  57.6,
  207,
  251.7,
  269.1,
  248.6,
  285.5,
  413.8,
  464.2,
  417.8,
  516.4,
  485.7,
  288.1,
  190.1,
  217.4,
  287.5,
  200,
  77.9,
  45.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.4,
  23.5,
  49.4,
  106,
  139,
  114.4,
  113.9,
  144.7,
  177.2,
  206.3,
  191.8,
  148,
  253.5,
  253.4,
  123.8,
  166.2,
  180.1,
  136.9,
  138.9,
  111.2,
  84.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.3,
  19.4,
  44.1,
  77.4,
  117,
  162.9,
  186,
  231.5,
  329.4,
  502.2,
  492.1,
  505.4,
  509.5,
  490.6,
  459.4,
  416.7,
  374.4,
  319.9,
  245.3,
  175.3,
  110.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  10.8,
  53.5,
  106.3,
  209,
  255.5,
  328.6,
  390.4,
  445.1,
  492.1,
  522.1,
  549.7,
  558.3,
  551.6,
  527.3,
  494.9,
  458.6,
  416.3,
  357.6,
  279.2,
  205.8,
  122.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.7,
  12.1,
  31.9,
  46,
  63,
  104,
  125.2,
  140.6,
  176.4,
  213.7,
  201.1,
  234,
  495.2,
  464.4,
  459.1,
  422.5,
  370.1,
  312.3,
  248,
  178.7,
  112.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.2,
  21.5,
  44.8,
  80.7,
  115.3,
  145.8,
  171.6,
  278.2,
  439,
  505.5,
  532.3,
  522.9,
  519.7,
  508.5,
  483.9,
  443.7,
  393.3,
  335.9,
  271.5,
  174.3,
  109.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  14.3,
  54.7,
  114.3,
  187.3,
  254.8,
  319.9,
  387.4,
  443.1,
  499.6,
  529.7,
  543.3,
  428.1,
  301.3,
  218.4,
  374.1,
  354.3,
  203.5,
  183,
  184.6,
  164.2,
  108.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.6,
  17,
  30.1,
  38.8,
  38,
  46.9,
  37.6,
  35.7,
  31,
  44.4,
  49.2,
  52.3,
  68,
  53.1,
  49.8,
  69.5,
  52.7,
  51.7,
  23.9,
  29.6,
  63,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.5,
  17.9,
  58,
  134.3,
  163.8,
  86.7,
  102.7,
  162.1,
  108.8,
  82.8,
  51,
  40.4,
  33.8,
  46.6,
  56.8,
  49.6,
  38.7,
  21,
  17,
  24.7,
  18.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.2,
  5.5,
  7,
  9,
  15.3,
  18.4,
  46.8,
  48.7,
  46,
  42.1,
  55.6,
  64.8,
  45.4,
  49.7,
  41.8,
  49.7,
  54.7,
  32.1,
  34.8,
  16,
  20.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.4,
  10.7,
  33.1,
  107.7,
  157.5,
  156.1,
  149.9,
  177,
  146.8,
  199.7,
  277.9,
  238.5,
  364.2,
  374.6,
  329.3,
  263.7,
  326.4,
  432.8,
  123,
  111.9,
  108.9,
  75.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.3,
  10,
  37.8,
  66.4,
  44.2,
  21.8,
  63.2,
  71.8,
  70.8,
  76.1,
  99.2,
  89.4,
  61,
  30.4,
  65.9,
  57.4,
  72.7,
  66.2,
  26.3,
  23.8,
  13.8,
  11.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.1,
  4.5,
  11.8,
  15.2,
  91.6,
  62.5,
  57,
  46.8,
  103.8,
  125.3,
  246.3,
  132.8,
  119.9,
  121.9,
  289.5,
  138.4,
  222.8,
  133.6,
  55.1,
  63.7,
  17.8,
  23,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.9,
  19.9,
  77.6,
  189.9,
  149.6,
  157.1,
  163.9,
  225.3,
  289.2,
  234.2,
  289.8,
  315.4,
  164.3,
  134,
  102.5,
  108,
  59,
  74.7,
  80,
  77.2,
  82.4,
  14.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.1,
  17.1,
  66.4,
  45,
  100,
  115.8,
  236.7,
  174.1,
  205,
  385.9,
  430.2,
  165.1,
  280.6,
  380,
  197.6,
  363.4,
  359,
  412.6,
  375.8,
  165.8,
  224.3,
  127.4,
  37.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  13.9,
  59,
  145.4,
  109.9,
  228,
  346.5,
  296.9,
  296.4,
  273.6,
  283.6,
  453.1,
  545.6,
  661.1,
  522,
  654.1,
  509.7,
  617.3,
  530.4,
  426.4,
  344.8,
  275.1,
  140.3,
  112.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.4,
  9.8,
  10.6,
  22.4,
  46.4,
  67.1,
  28.8,
  33.3,
  68.5,
  55.1,
  87.4,
  94.1,
  75.2,
  87.2,
  85.6,
  58.6,
  43.2,
  28.6,
  20.7,
  10.6,
  7.9,
  5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.2,
  19.9,
  41.2,
  51.5,
  50.6,
  46.5,
  73,
  143.4,
  114.5,
  176,
  143.7,
  116,
  178.6,
  96.8,
  131.2,
  138.5,
  134.6,
  106.8,
  73.2,
  59.7,
  52.6,
  19.8,
  7.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.3,
  19.1,
  16.4,
  22.9,
  61,
  138.3,
  235.9,
  240.9,
  106.8,
  146.4,
  219.8,
  228.2,
  131.3,
  222.9,
  202.1,
  213,
  161.5,
  195.4,
  164.9,
  106.4,
  86,
  62.5,
  49.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  9.4,
  36.5,
  62.5,
  117.1,
  142.5,
  175.1,
  197.2,
  249.7,
  331.8,
  197.5,
  138.7,
  144.3,
  180.6,
  185.2,
  181.2,
  145.8,
  150.9,
  137.3,
  115.5,
  78.7,
  80.7,
  34.1,
  32.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  14.8,
  51.9,
  100.8,
  154.9,
  260.4,
  360.4,
  403.8,
  356.7,
  562.7,
  456.1,
  386.5,
  369.5,
  551.2,
  461.7,
  396.3,
  562.7,
  470.7,
  428.7,
  327.7,
  390.8,
  235,
  155.3,
  49.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  13.2,
  20.8,
  72.4,
  90.3,
  83.9,
  192.9,
  206.1,
  340.9,
  259.1,
  350.3,
  384.8,
  398.5,
  288.6,
  385.3,
  198.8,
  207.7,
  220.5,
  216.2,
  237.9,
  192.6,
  129.6,
  67.6,
  39.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.6,
  23.6,
  60.1,
  78.6,
  113.7,
  132.8,
  215.1,
  319.5,
  370.3,
  423.1,
  384.7,
  299.9,
  445.9,
  302.9,
  305,
  279.5,
  115.6,
  70.5,
  153,
  98.7,
  113.9,
  101.4,
  52.8,
  45.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.5,
  35.8,
  99.6,
  162.2,
  231.7,
  317.8,
  421.4,
  488.7,
  376.5,
  399.8,
  547.1,
  656.5,
  581.6,
  638.7,
  341.9,
  191.7,
  360.1,
  631.1,
  338.2,
  424.1,
  421,
  333.1,
  253.8,
  172.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.5,
  30.9,
  87.8,
  158.3,
  226.1,
  304.1,
  386.5,
  457.4,
  515.5,
  566.3,
  615.1,
  642.6,
  658.2,
  659.7,
  616.9,
  641.8,
  585.2,
  558.6,
  480.7,
  457,
  387.1,
  311.4,
  235.5,
  156.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.3,
  36.1,
  89.9,
  159,
  235.9,
  308.9,
  388.5,
  462.7,
  525.8,
  578.1,
  622.6,
  648.4,
  666.9,
  662.4,
  651.3,
  634.2,
  593.9,
  557.2,
  511.7,
  438.3,
  377,
  316.3,
  239.1,
  159.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5,
  22.5,
  50,
  86.8,
  119.5,
  135.5,
  158.3,
  184,
  213.5,
  220,
  256,
  305.3,
  329.1,
  401,
  403.2,
  422.9,
  313.5,
  252.2,
  209.4,
  196.7,
  204.6,
  163.3,
  126.3,
  93.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.7,
  19.5,
  29.6,
  55.1,
  74.8,
  232,
  322.7,
  185,
  188.3,
  220,
  293.7,
  342.1,
  126.7,
  101.7,
  72.8,
  67.7,
  216.6,
  272.3,
  308.6,
  415.4,
  414.2,
  356.7,
  217.9,
  144.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.4,
  24.9,
  45.4,
  104.7,
  189.7,
  140.1,
  364.2,
  146.6,
  456.1,
  451.3,
  362.9,
  550.4,
  354.4,
  393.8,
  534.7,
  398.1,
  396.1,
  216.3,
  296.4,
  178.5,
  216,
  185.5,
  105.5,
  179.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.4,
  2.2,
  5.6,
  9.4,
  9.8,
  16.4,
  27.3,
  35.6,
  38,
  50.8,
  52,
  50.1,
  49,
  40.3,
  54.8,
  45.9,
  49,
  52.2,
  42.1,
  31.4,
  20.1,
  18.8,
  12.5,
  13.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  11.7,
  29.2,
  97.7,
  210.2,
  291.4,
  346.7,
  480.1,
  551.4,
  496.9,
  556.8,
  602.1,
  595.5,
  730,
  555.7,
  502.7,
  521.8,
  405.2,
  457.8,
  456.6,
  441.7,
  450.9,
  373.9,
  344.7,
  167.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  18.2,
  63,
  137.5,
  225.4,
  300.7,
  384.9,
  465.8,
  533.3,
  590.5,
  646.3,
  683.8,
  718,
  674,
  721,
  569.5,
  537.3,
  672.3,
  642.5,
  581.9,
  522.8,
  457,
  379.6,
  295.8,
  206.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  19.9,
  76.8,
  144.1,
  219.8,
  295.8,
  367.8,
  441.1,
  502.3,
  585.5,
  631.8,
  674.5,
  707,
  740,
  653.7,
  728,
  707,
  660,
  628.4,
  569.4,
  511.8,
  418.4,
  322.9,
  233.5,
  152.3,
  83.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  12.2,
  40.3,
  98.8,
  140,
  165.5,
  212.1,
  264.2,
  306.4,
  432.4,
  460.4,
  445.5,
  470.6,
  567.2,
  540.3,
  551.5,
  519.7,
  611.6,
  561.1,
  406.1,
  326.5,
  296.9,
  283.9,
  263.4,
  194.1,
  109.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  18.9,
  48,
  79,
  112,
  124.1,
  236.9,
  448.1,
  486.7,
  526.4,
  560.8,
  599.5,
  644.5,
  643.7,
  678.7,
  635.1,
  604.8,
  634.7,
  602,
  447.5,
  363.8,
  391.7,
  324.7,
  246.5,
  163.8,
  99,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.9,
  6.5,
  12.6,
  52.3,
  52.9,
  85.6,
  256.3,
  229.1,
  75,
  61.1,
  245.5,
  101,
  199.2,
  140.4,
  280.9,
  263.4,
  255.3,
  529.8,
  290.8,
  429.1,
  530.4,
  297,
  201,
  131.4,
  128.8,
  74,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.7,
  16.2,
  69.3,
  132,
  166.5,
  127.3,
  171.9,
  193.4,
  357.1,
  274.8,
  254.5,
  640.4,
  406.1,
  255.5,
  745,
  517.3,
  516.8,
  447.2,
  327.4,
  467.1,
  335.4,
  183.2,
  218.1,
  120.2,
  136.5,
  50.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.7,
  52.4,
  138.3,
  258.9,
  268.6,
  325.7,
  409.1,
  396.6,
  308.1,
  296.2,
  302.4,
  368.6,
  451,
  499.5,
  645.3,
  696,
  462.8,
  472.7,
  606.1,
  281.3,
  297.5,
  135.9,
  89.3,
  74.1,
  40.9,
  24.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.5,
  4.6,
  22.2,
  86.6,
  95,
  57.7,
  100.2,
  368.3,
  523.9,
  497.6,
  359.2,
  185.7,
  177.2,
  181.7,
  57.2,
  161,
  146,
  163.4,
  125,
  163.6,
  87.6,
  75.4,
  241,
  147.3,
  59.2,
  55.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.3,
  18.8,
  50.1,
  75,
  73,
  204,
  171.6,
  333.5,
  289.9,
  284.2,
  417,
  358.5,
  452.5,
  480.5,
  572.5,
  594.6,
  568.8,
  527.5,
  431.3,
  341.3,
  381.2,
  403.8,
  206.8,
  155.6,
  96.3,
  68.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.3,
  10.1,
  23.2,
  63.5,
  100.6,
  136.3,
  141.9,
  184.6,
  275.6,
  235.9,
  268.4,
  390.7,
  494.4,
  330.3,
  441.4,
  327.3,
  243.9,
  226.6,
  181.7,
  136.8,
  198,
  219.4,
  183.4,
  173.9,
  204.6,
  152.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.7,
  50.3,
  122.9,
  211.6,
  280.8,
  349.6,
  422.3,
  502.2,
  578.4,
  641.1,
  687.9,
  734,
  765,
  782,
  790,
  780,
  753,
  728,
  684.3,
  633.8,
  564.3,
  497.5,
  419.5,
  337.9,
  252.2,
  165.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.9,
  28.5,
  70.3,
  107.7,
  209.3,
  216.7,
  173.2,
  66.1,
  101.6,
  115.7,
  85.8,
  136.9,
  240.7,
  138.3,
  131.2,
  120.7,
  220,
  443.7,
  205.3,
  330.4,
  350.6,
  301.8,
  478.8,
  370.8,
  288.1,
  198.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.6,
  22.2,
  41.6,
  73.2,
  104.9,
  160.4,
  163.6,
  224.4,
  231.6,
  252.5,
  214.8,
  219.3,
  263.6,
  212.9,
  196.5,
  176.1,
  209.4,
  114,
  165.3,
  312.8,
  188.3,
  190.5,
  132,
  299.7,
  91.2,
  155.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  14.1,
  62.5,
  128.6,
  207.1,
  286.7,
  369.5,
  458.7,
  572.5,
  611.4,
  582.2,
  788,
  611.1,
  705,
  743,
  965,
  644.5,
  609.8,
  363.2,
  503.1,
  413,
  331.8,
  283.5,
  197.4,
  200.9,
  100.2,
  141.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  14.3,
  62.9,
  128.7,
  210.3,
  295.4,
  353.8,
  443.1,
  528.7,
  595.7,
  663.4,
  720,
  760,
  800,
  809,
  734,
  801,
  770,
  736,
  679.5,
  600.1,
  593.1,
  517.5,
  424.2,
  344.6,
  249.7,
  190.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  19.8,
  83.4,
  150.6,
  128.8,
  187.2,
  365,
  242.7,
  61.5,
  164.8,
  291,
  413,
  342.9,
  433.4,
  249.6,
  259.9,
  324.9,
  362.4,
  248.7,
  300.5,
  542,
  301.9,
  505.3,
  210.7,
  177.4,
  156.2,
  60.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.9,
  23.9,
  68.5,
  138.7,
  209.5,
  294.1,
  338.3,
  426,
  522.2,
  614.2,
  661.5,
  720,
  763,
  792,
  781,
  825,
  755,
  649.9,
  689,
  714,
  629.7,
  568.1,
  482.5,
  414.8,
  322.3,
  249.9,
  174.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  22.3,
  64.7,
  131.3,
  165.6,
  257,
  350.5,
  514.1,
  328.2,
  309,
  417.4,
  587.5,
  558.1,
  478.3,
  484.3,
  534.9,
  455.4,
  404.2,
  320.5,
  392.4,
  352.1,
  381.3,
  372.3,
  334.1,
  336.7,
  242.2,
  167.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.9,
  16.3,
  37.3,
  56.9,
  72.4,
  82.3,
  171.7,
  231.9,
  229.1,
  280.2,
  276.6,
  232.6,
  201.7,
  187.2,
  215.3,
  203.4,
  117.5,
  268.1,
  172.4,
  204.9,
  163.4,
  196.2,
  178,
  190.7,
  102.2,
  68.4,
  42,
  26.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  10.7,
  27.3,
  54.6,
  99.6,
  220,
  335.8,
  318,
  498.7,
  358.3,
  408.6,
  474,
  426.8,
  446.3,
  479,
  420.3,
  463.8,
  432.1,
  485.6,
  271.7,
  204.4,
  240.3,
  250,
  199.3,
  205.6,
  109,
  46.8,
  30.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  4.2,
  19.3,
  32.1,
  31,
  57.7,
  91.2,
  95.1,
  122.5,
  146.2,
  209.5,
  265,
  197,
  150.8,
  308.8,
  164.2,
  208.5,
  271.3,
  382.9,
  262.1,
  78.3,
  38.1,
  126.2,
  146.6,
  117.2,
  93.1,
  55,
  8.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.4,
  43.4,
  48.9,
  71.8,
  102,
  33.2,
  45.1,
  52.3,
  45.8,
  64.3,
  45.4,
  114.2,
  64.1,
  43.7,
  82.5,
  87.5,
  71.4,
  85.8,
  98.2,
  101.7,
  74.2,
  162.1,
  150.7,
  113.5,
  92.9,
  59.5,
  32.1,
  19.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.9,
  3.5,
  5,
  9.7,
  16.8,
  20.7,
  35.2,
  29.3,
  64.7,
  53.3,
  53.2,
  59.5,
  60.5,
  80.5,
  66.6,
  44.7,
  40.5,
  55.1,
  63.9,
  72.5,
  77,
  52.7,
  25.5,
  33,
  37.4,
  15.1,
  14.5,
  5.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.6,
  24.4,
  27.6,
  65.4,
  78.2,
  152.6,
  160.6,
  224.4,
  242.9,
  231.5,
  379.6,
  518.3,
  568.1,
  551.2,
  487,
  374.9,
  358.5,
  336.2,
  298.4,
  243.5,
  218,
  249.2,
  143.9,
  102.6,
  64.6,
  56.7,
  62.4,
  49.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.5,
  32.1,
  82.5,
  144.7,
  214.8,
  280.9,
  341.8,
  440.3,
  546.5,
  616.8,
  685.5,
  732,
  760,
  406.3,
  548.7,
  628.2,
  374.7,
  728,
  817,
  655.4,
  422.9,
  322.6,
  218.9,
  186.9,
  168.4,
  167.8,
  159.1,
  105.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6,
  36.5,
  74.6,
  184.1,
  261.7,
  333.9,
  374.2,
  457.1,
  517.2,
  596.2,
  641,
  732,
  770,
  807,
  803,
  810,
  802,
  779,
  734,
  688.6,
  633,
  565.5,
  492.6,
  421.6,
  334.6,
  251.3,
  172.2,
  100.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.7,
  39,
  89.6,
  143.6,
  191.2,
  221.2,
  359.6,
  423.6,
  510.8,
  515.8,
  587.1,
  589.8,
  682.3,
  732,
  753,
  746,
  719,
  695.2,
  650.8,
  663.7,
  559.8,
  500.5,
  394,
  363.5,
  266.3,
  188.6,
  120,
  73.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.9,
  49.1,
  52,
  75.2,
  95,
  60.9,
  73,
  85.9,
  89.1,
  177.9,
  356,
  453.1,
  349.5,
  261.3,
  684.3,
  324.7,
  168.9,
  181,
  62.8,
  87.9,
  96.3,
  92.2,
  47.9,
  59.9,
  54,
  32.6,
  35.9,
  67.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.8,
  14.9,
  37.2,
  45.5,
  54.5,
  72.5,
  48.2,
  35.1,
  186.3,
  195.5,
  241.9,
  192.1,
  279.8,
  197,
  104.3,
  645.2,
  205,
  55.6,
  66.8,
  152.6,
  132.3,
  263.8,
  327.7,
  270.2,
  234,
  175.3,
  83.9,
  109.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.5,
  3.3,
  9.2,
  9.4,
  27.2,
  40.8,
  54.3,
  52.9,
  42,
  43.6,
  75,
  112.6,
  109.8,
  92.2,
  106.4,
  65.5,
  104.5,
  123.7,
  195.5,
  172.3,
  177.1,
  182.3,
  188.9,
  156,
  203.9,
  167.7,
  168.6,
  133.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  13,
  58.8,
  119.1,
  197.8,
  273.8,
  369.1,
  420.4,
  429.6,
  326.1,
  460.2,
  478.3,
  167.6,
  519.4,
  309.4,
  333.7,
  345.8,
  153.6,
  309.8,
  240,
  298,
  416.2,
  665.6,
  514,
  208.7,
  387.5,
  322.2,
  219.1,
  198.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  13.4,
  58,
  113.2,
  160.8,
  261,
  396.9,
  433.6,
  378.2,
  358.3,
  382.3,
  366.1,
  440.6,
  256.3,
  148.8,
  108.4,
  93.9,
  267.1,
  358.5,
  300.1,
  241.4,
  273.8,
  180,
  265.1,
  110.8,
  63.3,
  235.1,
  176,
  93.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3,
  8.6,
  22.1,
  35.9,
  77,
  167,
  246.6,
  77.6,
  58.6,
  539.8,
  447.4,
  234.6,
  252.6,
  319.1,
  154.6,
  464.8,
  390.4,
  581,
  380.7,
  131.6,
  132.4,
  52.8,
  88.4,
  224.9,
  157.5,
  149.9,
  185.6,
  167.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  5.9,
  21.3,
  29.3,
  60,
  72.5,
  125.4,
  209,
  315.9,
  327.5,
  365.4,
  472.4,
  379.6,
  554.5,
  382.2,
  587.4,
  232.2,
  494.8,
  488.8,
  352.3,
  314.5,
  395.2,
  379,
  350.9,
  377.2,
  197.7,
  146.7,
  150,
  156.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  11.2,
  21.6,
  70.9,
  143.2,
  176.5,
  171.2,
  284.2,
  233.6,
  252.7,
  329.7,
  307.2,
  327.3,
  415.2,
  281.5,
  228.4,
  215.4,
  286.8,
  270.7,
  274,
  148.8,
  72.2,
  89.7,
  161.8,
  326.3,
  113.3,
  45.7,
  7.7,
  9.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  21,
  89.6,
  134.1,
  178.8,
  268.2,
  367.7,
  452.3,
  292.5,
  144.8,
  314,
  327.7,
  410.1,
  378.8,
  467.6,
  797,
  286.7,
  795,
  625,
  486.6,
  571.3,
  521.6,
  354.8,
  331.3,
  463.7,
  387.7,
  175.1,
  67.8,
  42.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.2,
  18.8,
  67.5,
  133.8,
  207.1,
  285.2,
  367.5,
  441.9,
  460.5,
  558.7,
  497.6,
  705,
  740,
  576.8,
  446,
  743,
  777,
  833,
  659.3,
  652.3,
  628.4,
  478.4,
  553.6,
  249.1,
  181.5,
  293.7,
  190.8,
  173.8,
  102.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.6,
  5.7,
  11.2,
  35.5,
  18.5,
  23.3,
  44.1,
  72.4,
  65.9,
  46.7,
  54.7,
  66.5,
  40.7,
  52.1,
  38.4,
  79.5,
  80.1,
  52.9,
  64.9,
  81.8,
  77.3,
  66.3,
  73.7,
  84,
  117.6,
  95.8,
  95.3,
  94.9,
  108.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.5,
  34.8,
  82.8,
  142.8,
  200.7,
  215.7,
  178.7,
  208.4,
  231.1,
  387,
  615.1,
  705,
  735,
  785,
  821,
  831,
  492.7,
  616.5,
  742,
  562.8,
  668.5,
  323.7,
  403.4,
  475.4,
  409.8,
  387.8,
  299.9,
  220.6,
  145.3,
  75.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.7,
  19.4,
  80.3,
  106.8,
  150.9,
  258.1,
  336.9,
  432.2,
  443.5,
  496.8,
  621.8,
  671.6,
  658.2,
  746,
  771,
  779,
  772,
  677.7,
  540.4,
  457.5,
  628.7,
  618.7,
  566.6,
  384.8,
  438.6,
  355.8,
  232.3,
  174.7,
  129.1,
  81.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.5,
  20.6,
  53.5,
  113,
  184.5,
  263.6,
  355.8,
  387.4,
  476.7,
  530.5,
  550.8,
  671.1,
  720,
  764,
  793,
  808,
  815,
  809,
  788,
  743,
  717,
  663.6,
  608.9,
  556.3,
  528.4,
  442.6,
  352.3,
  343.5,
  233.1,
  51.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.7,
  30.1,
  53.7,
  64.3,
  170.8,
  174.6,
  172.3,
  160.9,
  222.8,
  343.8,
  616.2,
  465.6,
  668,
  710,
  705,
  381.2,
  259.8,
  247.6,
  135.4,
  114.3,
  58.5,
  176,
  193.8,
  194.1,
  130.9,
  147.3,
  129.5,
  91.3,
  70.2,
  22.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2,
  14.4,
  32.6,
  78.2,
  134.1,
  202.3,
  213.6,
  344.5,
  276.2,
  192.9,
  451.5,
  599.8,
  481.8,
  613.3,
  677,
  752,
  548.1,
  620.9,
  753,
  728,
  802,
  591.3,
  560.2,
  589.2,
  464.6,
  429,
  349.2,
  195,
  184.6,
  75.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.6,
  18.4,
  36,
  73.5,
  125.7,
  158.6,
  240.5,
  320.3,
  423,
  407.3,
  481,
  556.1,
  344.7,
  371.3,
  600.2,
  940,
  818,
  564.2,
  256,
  10.4,
  52.2,
  120.5,
  145.7,
  118.8,
  84.9,
  98.2,
  63.8,
  94.3,
  43.5,
  9.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.2,
  32.2,
  29.1,
  18.4,
  38.7,
  58.7,
  62.3,
  88.6,
  152.3,
  182.3,
  136.4,
  167.7,
  160.8,
  181.9,
  325,
  315.2,
  305.2,
  822,
  705,
  363.8,
  127.4,
  341.7,
  122.6,
  94.1,
  42.8,
  42.9,
  102.8,
  99.6,
  29.2,
  9.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.7,
  4.9,
  13.3,
  47.6,
  90.2,
  91.3,
  128.9,
  51.1,
  224,
  227.8,
  149.4,
  201.2,
  214.6,
  174.4,
  215.6,
  459,
  171.9,
  216.4,
  203.1,
  116.6,
  169.9,
  265.3,
  146.8,
  153.8,
  97.6,
  90.2,
  74.3,
  117.4,
  45,
  36.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  9.9,
  45.6,
  103.4,
  178.4,
  244,
  334.9,
  471.1,
  326.7,
  173.5,
  234,
  374.5,
  565.4,
  363.4,
  281.6,
  723,
  567.7,
  829,
  529.5,
  352.4,
  435.1,
  291.2,
  429.9,
  214.1,
  442.5,
  379.2,
  409.6,
  382.4,
  298.6,
  214.6,
  137.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  14.6,
  63.2,
  155.9,
  170.4,
  218.1,
  287.9,
  310.8,
  503.3,
  222.1,
  451.9,
  222.6,
  451.4,
  407.1,
  555.8,
  440.5,
  599.1,
  752,
  746,
  749,
  735,
  666.2,
  542.3,
  681.9,
  508.6,
  484.5,
  498.1,
  277.7,
  312.4,
  85.5,
  111.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  8.9,
  38,
  105.9,
  176.8,
  238,
  334.7,
  363.7,
  475.1,
  591.4,
  585.6,
  664.8,
  488.6,
  509.9,
  783,
  619.3,
  637.1,
  747,
  838,
  862,
  832,
  760,
  748,
  679.7,
  555.8,
  523.7,
  394.6,
  357.2,
  240.6,
  222.1,
  126.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.2,
  11.1,
  47.9,
  121.3,
  183.4,
  165.8,
  230.7,
  234.9,
  294,
  311.9,
  319.3,
  338.3,
  395.3,
  471.4,
  682.9,
  672.2,
  694.6,
  838,
  680.8,
  562.9,
  436.5,
  445.7,
  404.6,
  370.6,
  261,
  227.9,
  191.4,
  135.2,
  67.6,
  44.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.9,
  6.4,
  20,
  15.5,
  32.4,
  64.6,
  49.3,
  76.8,
  86.6,
  109.1,
  169.4,
  155.4,
  165.8,
  129.2,
  215.5,
  142.2,
  178.8,
  185.6,
  189.3,
  185.1,
  148.3,
  135.5,
  175,
  187.2,
  210.3,
  153.1,
  153.1,
  90.7,
  52.9,
  34.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.8,
  26.2,
  46.6,
  77.1,
  100.9,
  128.1,
  194.8,
  376.1,
  392.7,
  542.6,
  374.3,
  267.3,
  302.8,
  390.1,
  397.6,
  499.8,
  563.3,
  442.1,
  367.9,
  401.1,
  347,
  469.4,
  692.8,
  683.5,
  363.8,
  390.8,
  395.3,
  302.4,
  215.2,
  132.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.8,
  24.9,
  64.9,
  118,
  181.9,
  214.3,
  223.7,
  277.2,
  370,
  382.8,
  553.6,
  747,
  788,
  814,
  802,
  797,
  829,
  850,
  815,
  743,
  757,
  719,
  681.1,
  598.4,
  535.7,
  444,
  369.1,
  289.8,
  221.3,
  150.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  8.1,
  26.1,
  65.1,
  152.9,
  244.3,
  245.9,
  411.8,
  511.1,
  585.1,
  648.5,
  717,
  771,
  819,
  856,
  887,
  895,
  901,
  893,
  880,
  850,
  801,
  748,
  687.7,
  617.4,
  548,
  466.3,
  385.3,
  298.9,
  221.6,
  145.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  9.2,
  29.3,
  86.3,
  176.1,
  181.6,
  304.4,
  436.3,
  503.5,
  582.6,
  651.6,
  713,
  769,
  805,
  842,
  877,
  867,
  861,
  901,
  872,
  775,
  769,
  727,
  574.3,
  619.7,
  551.1,
  486.9,
  322.4,
  228.7,
  152.4,
  121.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  17,
  57.3,
  114.3,
  186.9,
  263.7,
  348.4,
  429.1,
  512.7,
  590.8,
  695.7,
  666.7,
  806,
  792,
  792,
  797,
  870,
  820,
  737,
  868,
  767,
  800,
  565.2,
  592.4,
  308.9,
  372.9,
  252.7,
  226.8,
  89.2,
  150.1,
  38.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  15.2,
  51.5,
  104,
  176.9,
  256.7,
  336.2,
  418.5,
  497.8,
  573,
  642.4,
  704,
  763,
  786,
  854,
  863,
  875,
  880,
  819,
  887,
  850,
  811,
  748,
  680.4,
  617.8,
  546.5,
  469.7,
  390.1,
  305.7,
  224.9,
  151.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  17.1,
  57,
  110.6,
  185,
  265.8,
  346.4,
  428.2,
  509.8,
  586.1,
  654.7,
  718,
  781,
  827,
  865,
  889,
  906,
  907,
  899,
  878,
  842,
  804,
  753,
  690.2,
  625.2,
  553.1,
  472.4,
  392.4,
  232.9,
  186.6,
  150.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.1,
  15.4,
  55.2,
  107.5,
  180.3,
  258.4,
  338.1,
  416.1,
  492.5,
  563,
  623.8,
  701,
  730,
  668.5,
  448.8,
  253.2,
  258.5,
  457.9,
  429.2,
  491.3,
  573.4,
  268.3,
  420.9,
  533.8,
  398.2,
  216.7,
  200.6,
  335.8,
  289.9,
  186.5,
  125.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.3,
  20.5,
  56.3,
  97.2,
  146.4,
  224.4,
  312.1,
  397.1,
  494.4,
  555,
  592.8,
  595.9,
  699.3,
  691.6,
  507.3,
  935,
  935,
  902,
  850,
  823,
  773,
  764,
  729,
  483.8,
  647.7,
  482.2,
  382,
  304.6,
  157.3,
  134.5,
  82.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3,
  27.5,
  60.5,
  142.5,
  116.4,
  227.2,
  265.8,
  187.9,
  334.9,
  335.9,
  440.7,
  514.2,
  741,
  790,
  717,
  810,
  802,
  776,
  800,
  724,
  731,
  604.9,
  463.4,
  597.3,
  562.8,
  256.4,
  235.2,
  236.4,
  186.4,
  183.5,
  147.8,
  67.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  15.1,
  67.1,
  114.2,
  68.7,
  161.1,
  330.8,
  406.5,
  493.5,
  578.3,
  624.3,
  680,
  742,
  783,
  818,
  658.1,
  644.6,
  736,
  774,
  746,
  436,
  322.9,
  278.4,
  17.5,
  16.5,
  48.6,
  284.2,
  183.3,
  85.6,
  61.3,
  29.8,
  32.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.7,
  30.3,
  20.1,
  27.6,
  26.7,
  43.3,
  74.9,
  82.9,
  146.1,
  134.5,
  107.8,
  96.8,
  179,
  164.7,
  187,
  154.2,
  47,
  86.5,
  60.2,
  96.1,
  209.3,
  314.1,
  370,
  339.1,
  331.7,
  245.6,
  445.8,
  137,
  131.8,
  142.2,
  76.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.2,
  21.3,
  61.3,
  108.7,
  182.2,
  156.9,
  176.2,
  263.5,
  303.6,
  255.4,
  249.9,
  439.4,
  594.3,
  596.6,
  614.1,
  342.8,
  704,
  768,
  775,
  945,
  668.2,
  824,
  779,
  726,
  420.8,
  367,
  409,
  333.7,
  292.9,
  214.5,
  148.8,
  89.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.2,
  18.9,
  56,
  110.7,
  178.5,
  251.4,
  330.3,
  404.3,
  477,
  548.1,
  620.9,
  676.2,
  738,
  784,
  813,
  821,
  861,
  867,
  812,
  666.7,
  590,
  640.2,
  626.2,
  578,
  581.1,
  480.6,
  413.6,
  362.1,
  203.2,
  123.6,
  87.1,
  71,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.4,
  24.8,
  72,
  110.1,
  162.2,
  227.2,
  151.1,
  225.8,
  214.3,
  275.6,
  292,
  617.2,
  530.2,
  519.8,
  332.3,
  245.7,
  162.6,
  145.9,
  139.6,
  138.8,
  229.3,
  43.1,
  54.6,
  108.3,
  67.9,
  46.8,
  56.5,
  93.8,
  67.7,
  92.7,
  62.7,
  34,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  7.6,
  23.1,
  70.5,
  93.3,
  112.3,
  204.8,
  295.1,
  435.2,
  337,
  352.1,
  430.2,
  580.7,
  664.2,
  529.2,
  466.4,
  424.8,
  536.5,
  168.5,
  173.5,
  541.6,
  460.9,
  403.2,
  309.3,
  372.7,
  416.9,
  253,
  232.3,
  171.7,
  142.9,
  180,
  93.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  6.5,
  8.3,
  14.7,
  33.7,
  163.4,
  141.5,
  359.8,
  457.9,
  241.9,
  482.4,
  533.5,
  414.2,
  540.1,
  462.3,
  319.4,
  448.4,
  605,
  590.4,
  551.1,
  426.8,
  302.2,
  393.1,
  370.3,
  28,
  36.6,
  115.6,
  380.3,
  191.7,
  157.7,
  101,
  50.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  8.7,
  23.8,
  40.6,
  42.2,
  148.5,
  238.2,
  244.1,
  158.9,
  202.7,
  241.6,
  240.9,
  304.7,
  233.8,
  441.1,
  346.1,
  433.2,
  385.9,
  89.4,
  485,
  181.6,
  222.3,
  93.3,
  201.5,
  122.1,
  48.5,
  147.9,
  156.4,
  43.4,
  66.7,
  64.3,
  93.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.7,
  13.6,
  13.1,
  28.5,
  72,
  137.8,
  174,
  149.7,
  236,
  180.6,
  173.1,
  223.2,
  256.8,
  319.9,
  489.5,
  624.2,
  473.1,
  526.7,
  445.8,
  490.3,
  490.1,
  642.9,
  609.2,
  480.4,
  512.5,
  432.7,
  211.4,
  177.9,
  230.5,
  175.6,
  107.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.3,
  15.4,
  60.1,
  121.7,
  207,
  280.5,
  354.3,
  440.7,
  515.7,
  457.6,
  591,
  530.2,
  776,
  837,
  708,
  740,
  749,
  542.5,
  550,
  570.5,
  486.7,
  510.5,
  422.5,
  279.6,
  384.5,
  293.7,
  347.8,
  240.8,
  279.3,
  239.9,
  163.9,
  92.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.8,
  24.1,
  69.1,
  127.8,
  199.5,
  276.1,
  320,
  428.6,
  553.3,
  469.6,
  622.5,
  434.5,
  579.4,
  555.6,
  768,
  878,
  792,
  701,
  716,
  519.3,
  837,
  693.5,
  559.2,
  562,
  582.7,
  494.4,
  614.3,
  470.6,
  310.8,
  259.2,
  169.6,
  96.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6,
  22.9,
  29.8,
  32.3,
  46.9,
  49.3,
  63.7,
  229.6,
  468.1,
  487.4,
  502,
  356.6,
  279.1,
  493.3,
  545,
  329.5,
  452.5,
  560.9,
  766,
  317.8,
  315.5,
  653.2,
  624.1,
  829,
  371.9,
  406.9,
  456,
  420,
  326,
  194,
  133,
  52.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  20,
  60.3,
  83.4,
  172.8,
  222.5,
  312.5,
  398.5,
  442,
  499.2,
  554,
  681,
  715,
  737,
  727,
  819,
  592,
  611.8,
  599.4,
  680.8,
  673.9,
  641,
  606.1,
  367.1,
  454.5,
  361.1,
  302.9,
  285.1,
  208.5,
  143.5,
  102.8,
  55.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.3,
  20.9,
  48.1,
  30.7,
  23.4,
  82.1,
  94.1,
  175.9,
  152.3,
  342.7,
  409.2,
  560.4,
  427.3,
  401,
  768,
  550.8,
  508.4,
  472.9,
  215.7,
  526.6,
  557.9,
  514.1,
  430.4,
  565.8,
  244.6,
  177.2,
  80.1,
  111.8,
  142.3,
  38.8,
  16.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1,
  14.4,
  66.9,
  36,
  134.8,
  175.2,
  168.7,
  257.6,
  362,
  272.5,
  361.8,
  274.7,
  678.1,
  788,
  622,
  294.8,
  166.6,
  740,
  762,
  432.9,
  291.6,
  234.8,
  749,
  621.3,
  305.9,
  412.8,
  423.4,
  214.7,
  84.6,
  157.5,
  105.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.5,
  13.9,
  42,
  111.7,
  159.2,
  155.9,
  184.4,
  238.6,
  519.1,
  497.1,
  564.8,
  528.8,
  468.4,
  415,
  232,
  353.8,
  520.4,
  203.2,
  244,
  374.2,
  269.7,
  472.5,
  314.5,
  376.1,
  57.1,
  193.2,
  224.3,
  262,
  232.3,
  54.7,
  37.1,
  158.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.1,
  11.9,
  22.1,
  35.9,
  67.3,
  117.1,
  117.8,
  205.4,
  182.3,
  229,
  134.3,
  165.6,
  70,
  192.8,
  222.1,
  183,
  175.4,
  89.9,
  96.3,
  128.4,
  190.9,
  97,
  115.5,
  115.9,
  108.6,
  54.4,
  75.6,
  129.8,
  62.9,
  70.6,
  32.1,
  20,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  4.5,
  30,
  42.7,
  32.9,
  63.3,
  184,
  156.3,
  253.1,
  301,
  339.3,
  381,
  422.3,
  401.9,
  273.3,
  223.9,
  289.3,
  286.6,
  216.2,
  437.9,
  421,
  216.2,
  444.1,
  356.8,
  366.3,
  334.5,
  266.9,
  189.5,
  148.6,
  106.1,
  77.7,
  29.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.3,
  14.2,
  37,
  73.9,
  135.4,
  185.8,
  339.2,
  339.2,
  402.4,
  482.8,
  628.1,
  698.8,
  749,
  737,
  803,
  893,
  632.6,
  603.2,
  438.5,
  329.6,
  225.9,
  180,
  154.3,
  141.1,
  119.6,
  25.3,
  25.1,
  42.3,
  56.9,
  29.1,
  13.7,
  16.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.9,
  7.3,
  20.1,
  25.2,
  31.8,
  61.7,
  135.8,
  127.8,
  137.2,
  60.3,
  107,
  130.4,
  92.4,
  196.8,
  145.6,
  191,
  557.4,
  366.2,
  173.2,
  94.2,
  95.1,
  84.7,
  128.9,
  225.8,
  142.5,
  140.2,
  290.1,
  264.1,
  170.6,
  55.2,
  30,
  33.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.1,
  3.3,
  11.7,
  41.8,
  76.8,
  115.8,
  108.3,
  124.9,
  199.6,
  195.1,
  231.6,
  347,
  468.9,
  455.9,
  637.2,
  819,
  795,
  460.9,
  423.5,
  268.6,
  132.5,
  79,
  50.2,
  36.5,
  173.5,
  202.3,
  155.5,
  356.9,
  210.9,
  169.5,
  110.4,
  23.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.2,
  14.3,
  66.6,
  77.2,
  172,
  258.8,
  342.2,
  365,
  195.8,
  278.9,
  300.5,
  253.8,
  404.1,
  156.8,
  823,
  643.8,
  310.3,
  333.8,
  325.9,
  485.7,
  340.1,
  278.4,
  359.8,
  387.1,
  394,
  384.3,
  124.6,
  251.7,
  236.6,
  283.7,
  142.4,
  47.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  18.7,
  61.1,
  117.1,
  172.5,
  148.6,
  157.2,
  208.4,
  202,
  250.1,
  373.9,
  501.4,
  607.6,
  406.7,
  461.3,
  327.8,
  148.2,
  24,
  15.6,
  40.1,
  37.6,
  85.7,
  54.7,
  80.8,
  95.3,
  115.5,
  61.8,
  17.4,
  23.9,
  21.9,
  9.9,
  9.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.6,
  13.4,
  15.2,
  54.7,
  30.7,
  59.9,
  166.3,
  66.6,
  172,
  132.7,
  231.4,
  217.6,
  125.8,
  108.6,
  127.9,
  94.1,
  113.9,
  151.9,
  131,
  67.6,
  129.5,
  93.7,
  178.6,
  57.5,
  48.5,
  79.1,
  93.1,
  47.1,
  26.6,
  10.4,
  12.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2,
  25.4,
  32,
  27.5,
  82.6,
  107.5,
  186.3,
  209.2,
  246.4,
  231.2,
  373.9,
  214,
  193,
  143.1,
  230.8,
  225.4,
  730,
  479.3,
  611.6,
  695,
  718,
  711,
  706,
  630.1,
  414.6,
  30.5,
  268.8,
  196,
  334.8,
  186.1,
  17.5,
  14.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  10.7,
  75.2,
  104.4,
  121.1,
  123.1,
  282.7,
  341.3,
  442.5,
  449.8,
  410.7,
  502.5,
  639.9,
  830,
  718,
  787,
  727,
  747,
  710,
  441.9,
  303.4,
  155.8,
  95.4,
  100.1,
  64,
  54.1,
  49.3,
  32.3,
  36.2,
  24.8,
  24,
  11.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  11.6,
  58.1,
  146.5,
  155.8,
  182.5,
  265.6,
  359.7,
  470.9,
  518.4,
  582.3,
  608.5,
  454.3,
  759,
  611.3,
  497.5,
  830,
  765,
  550.7,
  406.3,
  377,
  381.7,
  499.9,
  375.1,
  325,
  287.9,
  244.6,
  289.1,
  142.4,
  64.3,
  20.5,
  26.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  17.8,
  44.6,
  85,
  142.5,
  243,
  232.7,
  241.1,
  300.7,
  296.8,
  545.8,
  642.6,
  677.9,
  612.2,
  699.5,
  630.4,
  676.7,
  212.7,
  194.6,
  768,
  736,
  810,
  564,
  699,
  397.2,
  562,
  156.9,
  90.1,
  92.4,
  97.6,
  83.1,
  37.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.5,
  21.4,
  55,
  92,
  100.3,
  96.8,
  140.6,
  226,
  287.2,
  309.3,
  402,
  652.5,
  205,
  191.6,
  277.9,
  193,
  34.8,
  77.6,
  180,
  158.3,
  65.6,
  52.1,
  46.8,
  101.8,
  156.1,
  245.3,
  222.6,
  287.6,
  218.7,
  132.3,
  114.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.1,
  3,
  20.8,
  56.5,
  104.7,
  217.7,
  346.6,
  406.5,
  403,
  360.6,
  500.2,
  428.8,
  331.3,
  306.3,
  180.2,
  189.5,
  283.7,
  293.9,
  158.2,
  392,
  221,
  129.8,
  92.7,
  69.4,
  64.6,
  177.8,
  133,
  115.1,
  51.2,
  90.2,
  70.5,
  23.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  5.9,
  14.6,
  27.5,
  30.4,
  32.7,
  37.3,
  74.6,
  254.1,
  354.5,
  504.4,
  426.8,
  644.4,
  610.2,
  816,
  496.1,
  468.2,
  481,
  361.6,
  419.6,
  436.7,
  540.2,
  376.1,
  419.5,
  392.7,
  405.3,
  488,
  413.1,
  332,
  254.6,
  177.2,
  106.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  6.1,
  13,
  34.8,
  54.5,
  83.4,
  102.8,
  131.3,
  128.4,
  143.1,
  149.7,
  140.1,
  174.2,
  187.4,
  272.3,
  334.1,
  457.3,
  524,
  623.4,
  415.9,
  484.2,
  594,
  393.5,
  399.4,
  359.2,
  368.5,
  363.5,
  437.6,
  209.6,
  230,
  153.4,
  109.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.3,
  4.8,
  11,
  24.9,
  38.7,
  50.6,
  85.1,
  140.4,
  138.2,
  131.3,
  190.5,
  204.1,
  181.7,
  221.1,
  293.8,
  351.2,
  385.2,
  294.5,
  394.8,
  264.6,
  406.2,
  523.3,
  459.9,
  527.5,
  418.9,
  404.2,
  407.3,
  393,
  234.4,
  176.9,
  117.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  8.8,
  33.8,
  49.4,
  69,
  83.7,
  100.7,
  137.9,
  157.5,
  244.7,
  582.2,
  682.6,
  732,
  772,
  716,
  634.6,
  922,
  743,
  723,
  686.4,
  745,
  390,
  403.1,
  570,
  280.1,
  469.5,
  477.9,
  349.3,
  257.8,
  102.2,
  149.1,
  74.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  11.3,
  50.3,
  113.3,
  162,
  234,
  314.9,
  393,
  471,
  545.4,
  607.7,
  671.2,
  732,
  788,
  809,
  744,
  816,
  625.6,
  878,
  890,
  626.9,
  686.1,
  631.7,
  211.5,
  536.3,
  401.4,
  164.9,
  334.7,
  308.6,
  222.1,
  131.2,
  74.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.5,
  8.5,
  20,
  22.9,
  37.4,
  48.7,
  73,
  178.5,
  252.4,
  249.9,
  466.5,
  627.6,
  765,
  672.2,
  770,
  654,
  938,
  656.9,
  788,
  324,
  139.5,
  145.6,
  230.2,
  359.9,
  543,
  433.9,
  340.3,
  255.7,
  183,
  102.7,
  72.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  7.7,
  33,
  62.8,
  125.3,
  174.6,
  227.8,
  331.1,
  402.6,
  324.9,
  504.7,
  444.2,
  582.2,
  577.6,
  334.8,
  288.1,
  548.5,
  655.3,
  466.6,
  585.4,
  624.1,
  598.8,
  638,
  525.4,
  432.5,
  157.2,
  88.1,
  53.2,
  62.9,
  1.8,
  15.5,
  40.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.8,
  27.3,
  80.1,
  102.6,
  164.6,
  238.6,
  339.5,
  400.3,
  418.4,
  577.3,
  398.9,
  198.3,
  421.6,
  541.5,
  600.1,
  869,
  885,
  555.9,
  610.6,
  498.6,
  453.5,
  253.4,
  517.9,
  405.5,
  378.9,
  240.2,
  204,
  250.6,
  214.3,
  145,
  67.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.1,
  18.8,
  41.8,
  64.1,
  55.5,
  148.6,
  233,
  195.2,
  281.3,
  418.2,
  461.3,
  488.3,
  266.1,
  234.3,
  444.7,
  281.6,
  288.2,
  302,
  483.5,
  678.7,
  846,
  674.6,
  364.6,
  43.1,
  23,
  34.7,
  69.9,
  162.2,
  177.1,
  87.4,
  47.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  10.5,
  33.3,
  55.5,
  113.5,
  164.5,
  248,
  191.8,
  81,
  98.3,
  87.6,
  164,
  367.7,
  393.3,
  165.6,
  259.3,
  338,
  386.6,
  324,
  441.9,
  384.6,
  540.5,
  293.5,
  284.2,
  275.4,
  261.9,
  187.6,
  164.7,
  176,
  61.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.1,
  22.7,
  49.9,
  70.6,
  138,
  226.8,
  236.6,
  369,
  379.2,
  482.7,
  278,
  389.2,
  357.4,
  246.4,
  388.2,
  652.8,
  317.2,
  194.5,
  314.8,
  388.9,
  125.4,
  163,
  158.9,
  82.9,
  47.3,
  46.1,
  92,
  72.2,
  64.9,
  47.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.4,
  16.3,
  33.4,
  46.6,
  108.4,
  156.1,
  148.5,
  158.2,
  104.9,
  278.4,
  381,
  383.4,
  510.4,
  563,
  593,
  394.7,
  283.5,
  93.9,
  326.3,
  170.2,
  360.8,
  184.5,
  158.1,
  96.6,
  116.7,
  219.9,
  59.3,
  122,
  36.7,
  36.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.2,
  22.7,
  43.1,
  99.6,
  153.2,
  250.8,
  315.8,
  381.7,
  485.7,
  579.6,
  617.3,
  601.7,
  786,
  731,
  601.3,
  778,
  310.1,
  114.6,
  512,
  471.1,
  525.3,
  375.3,
  499.8,
  483.8,
  437.8,
  419.2,
  339.4,
  353.6,
  199.3,
  139.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.8,
  15.7,
  39.3,
  85.8,
  134.2,
  142.6,
  214.3,
  328.5,
  373.7,
  437.4,
  721,
  786,
  640,
  696.6,
  880,
  536.5,
  267.3,
  232.4,
  115.2,
  376.5,
  476.8,
  76.9,
  137.1,
  418.4,
  92.2,
  186.7,
  169.3,
  246.5,
  142.9,
  162.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.7,
  11.6,
  44,
  59,
  56,
  76.9,
  181.8,
  368.4,
  459.9,
  352.5,
  370.7,
  472.9,
  529.9,
  440.3,
  405.3,
  340.1,
  414.3,
  362,
  222.6,
  141,
  98.6,
  113.9,
  148,
  96.7,
  161.2,
  112,
  72.3,
  86.7,
  29.8,
  21.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.1,
  14.9,
  30.5,
  51.5,
  50.9,
  86.8,
  153.9,
  151.3,
  165,
  302.2,
  270.9,
  357.6,
  346.1,
  519.1,
  549.4,
  488.1,
  565,
  294.1,
  147.9,
  73.6,
  173.2,
  308.2,
  413.5,
  88.2,
  392.1,
  443.6,
  255.9,
  221.9,
  85.5,
  96.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.8,
  25.1,
  81.3,
  117.7,
  184.1,
  276.1,
  346.8,
  451.2,
  357.7,
  490.6,
  477,
  634.7,
  682.4,
  599.5,
  764,
  753,
  670.7,
  684.4,
  699.1,
  777,
  682,
  638.3,
  665.5,
  589,
  527.1,
  397.4,
  364.1,
  274.6,
  196,
  114.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3,
  19.9,
  58.7,
  107.2,
  200.6,
  269.2,
  260.9,
  235.8,
  258.5,
  249.3,
  271.8,
  291.8,
  293.5,
  295.8,
  325.6,
  237.8,
  164.3,
  138.9,
  194.9,
  178.2,
  191.6,
  166.1,
  277.5,
  279.9,
  278.4,
  364.5,
  246.9,
  161.5,
  107.2,
  64.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.2,
  3,
  14.2,
  17.2,
  20.8,
  24.6,
  72.4,
  136.3,
  61.2,
  33,
  97.4,
  118,
  406.3,
  528.7,
  320.1,
  184.4,
  549.7,
  117.3,
  409.8,
  613.2,
  436.2,
  358.5,
  278.9,
  165.9,
  87.3,
  53.2,
  114.7,
  147.6,
  125.7,
  77.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.1,
  34.2,
  91.6,
  177.4,
  174.2,
  298.1,
  456.6,
  451.9,
  542.5,
  591.7,
  709,
  635.2,
  805,
  513.4,
  782,
  724,
  879,
  710,
  429.2,
  677.2,
  496.1,
  462,
  391.2,
  315.3,
  279.6,
  169.7,
  58.8,
  16.1,
  7.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.2,
  12.6,
  22.4,
  52.7,
  60.1,
  73.7,
  182.9,
  138.2,
  311.9,
  208.6,
  203.4,
  374,
  277.3,
  428.4,
  362.3,
  231.3,
  265.3,
  258.8,
  209.2,
  351.6,
  429.1,
  428.1,
  238.5,
  326.2,
  311,
  307.3,
  283,
  223.5,
  125.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.2,
  19.7,
  39,
  86.8,
  147.4,
  240.6,
  338.3,
  400.1,
  485.6,
  553.8,
  615.5,
  686.7,
  730,
  700,
  762,
  576.9,
  583.6,
  660.7,
  624.6,
  478.8,
  307.2,
  221.9,
  305.4,
  223.5,
  281.7,
  299.4,
  275.1,
  244.2,
  174.7,
  99.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  16.9,
  75.1,
  122.3,
  175.3,
  256.1,
  334.7,
  413.2,
  492.6,
  570.1,
  609.6,
  678.6,
  701,
  579,
  732,
  778,
  867,
  675,
  784,
  833,
  734,
  647.1,
  522.8,
  457.3,
  492.8,
  297.6,
  312.5,
  191.5,
  148.7,
  76.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2,
  18.5,
  57.1,
  124.1,
  122.6,
  246.2,
  325.9,
  332.6,
  315.8,
  339.6,
  347,
  522.9,
  642.9,
  380.3,
  372.8,
  395.8,
  299.7,
  248.6,
  109.6,
  122.8,
  87.9,
  45,
  88.6,
  169.3,
  203.9,
  359.7,
  230.2,
  208.4,
  219.5,
  144.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2,
  14.5,
  32.5,
  32.2,
  120.2,
  207.3,
  406.4,
  279.6,
  48,
  240.9,
  345.4,
  425.3,
  271.3,
  437.3,
  586,
  445.3,
  479.8,
  311.8,
  245.4,
  126.5,
  328,
  187.4,
  184.5,
  122.8,
  144.3,
  149.7,
  71.5,
  131.8,
  43.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.6,
  6.6,
  8.8,
  13,
  34.2,
  50.3,
  125.6,
  103.9,
  144.1,
  170.5,
  388,
  516.2,
  702,
  396.5,
  431.3,
  597.7,
  602.3,
  383.1,
  504.7,
  355,
  330.2,
  312.3,
  169.9,
  118.2,
  60.5,
  65.6,
  59.9,
  44.6,
  20.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.2,
  10.6,
  21,
  43.5,
  72.6,
  55,
  164.4,
  223.7,
  366.2,
  556.7,
  462.8,
  574,
  405.9,
  585.4,
  713,
  654.5,
  593.5,
  680.9,
  585.8,
  718,
  489,
  472.6,
  373,
  424.9,
  298.2,
  300,
  260.8,
  99.1,
  47.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  12.7,
  32.3,
  69.8,
  125.1,
  173.4,
  200.7,
  240.8,
  445.2,
  363.7,
  400.5,
  490.7,
  390.6,
  380.3,
  370.4,
  310.6,
  505.6,
  681.4,
  446.4,
  225.8,
  236.4,
  192.5,
  115,
  121.3,
  80.5,
  76.4,
  53.8,
  22,
  17.3,
  13.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.7,
  25.1,
  68.1,
  156.2,
  243.3,
  204.6,
  304.2,
  401.5,
  468.3,
  596.7,
  637.8,
  581.7,
  696.2,
  789,
  810,
  819,
  801,
  727,
  400.5,
  309.4,
  253.8,
  266.1,
  273.6,
  270,
  346.9,
  271.7,
  196,
  157.7,
  81.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  13.3,
  66.5,
  104.8,
  120.2,
  247.9,
  224.8,
  298.9,
  460.9,
  435.5,
  618.4,
  649.3,
  679.7,
  833,
  838,
  848,
  830,
  823,
  779,
  705,
  642.7,
  735,
  517.6,
  428.7,
  546.5,
  425.2,
  328,
  253.3,
  154,
  117.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.5,
  38.8,
  94.2,
  165.3,
  243.6,
  324.8,
  404.4,
  480.8,
  553.3,
  618.7,
  675,
  721,
  766,
  805,
  822,
  836,
  809,
  793,
  767,
  771,
  684.3,
  547.7,
  468.3,
  476.6,
  403.6,
  317.6,
  242.1,
  162.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.7,
  36.5,
  87,
  155,
  232.1,
  311,
  388.2,
  465.6,
  538.9,
  606.6,
  660,
  704,
  756,
  787,
  816,
  795,
  803,
  771,
  669.7,
  700,
  681.8,
  447.9,
  537,
  444.9,
  345.1,
  212.8,
  228.8,
  152.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.2,
  28.8,
  80.6,
  141.5,
  219.7,
  299.9,
  379.8,
  456.8,
  528.8,
  594.7,
  651.1,
  705,
  745,
  772,
  768,
  812,
  794,
  654.7,
  474.6,
  620.1,
  604.1,
  428.8,
  423.9,
  423.2,
  134.5,
  295.4,
  194.9,
  115.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.3,
  30.4,
  78.9,
  142,
  217.5,
  296.5,
  376.3,
  452.2,
  524.2,
  586.2,
  629,
  693.7,
  735,
  369.9,
  280.7,
  208.8,
  212.3,
  197.7,
  527.8,
  711,
  516.2,
  428.3,
  227.7,
  101,
  160.6,
  162.1,
  112.8,
  100.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.6,
  28.4,
  70.6,
  137.5,
  194.6,
  267.1,
  340.2,
  431.2,
  504.3,
  574.2,
  635.3,
  680.3,
  718,
  745,
  760,
  793,
  692.3,
  698.4,
  768,
  628.5,
  537.3,
  521.8,
  517.9,
  413.4,
  344,
  285,
  205.6,
  131.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.5,
  28.8,
  80.1,
  149.2,
  204,
  283.3,
  370.1,
  444.4,
  506.7,
  573.8,
  641.8,
  699,
  748,
  775,
  790,
  792,
  788,
  766,
  738,
  702,
  655.4,
  602.6,
  531.3,
  461.4,
  383.3,
  302.2,
  219.7,
  141.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.4,
  25.9,
  78.3,
  144.6,
  228.2,
  314.8,
  399.2,
  466.7,
  514.2,
  570.8,
  626.3,
  615.4,
  693.4,
  753,
  715,
  744,
  679.7,
  691.8,
  758,
  618.7,
  619.1,
  451.1,
  366.6,
  190.8,
  228.1,
  308.9,
  252.3,
  162.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.8,
  22.2,
  63.5,
  129.9,
  202.1,
  300.2,
  322.8,
  396.3,
  494.9,
  555.8,
  617.4,
  671.4,
  705,
  735,
  758,
  780,
  696.4,
  714,
  728,
  644.4,
  517.4,
  456.4,
  462.1,
  361.5,
  308.2,
  196.9,
  150.9,
  109,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.7,
  18.4,
  37.6,
  58.8,
  53.2,
  80.2,
  101.6,
  96.5,
  93.7,
  262.3,
  386.1,
  321.1,
  236.8,
  234.6,
  185.4,
  235.4,
  260.9,
  141,
  239.1,
  169.4,
  140.8,
  132.8,
  249.1,
  311.2,
  331,
  221.9,
  180.8,
  84.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.9,
  10.2,
  32.4,
  83.6,
  172.1,
  248,
  296.3,
  316.5,
  285.9,
  325,
  521,
  656.2,
  573.6,
  626.6,
  578.4,
  662.5,
  656.7,
  554.2,
  478.7,
  511.8,
  547.6,
  429.4,
  512.3,
  362.4,
  345.7,
  252.7,
  172.1,
  113.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.4,
  18.2,
  54.7,
  89.9,
  132.2,
  275.4,
  310.2,
  258.6,
  477.4,
  562.5,
  537,
  619.1,
  527.5,
  571.5,
  742,
  673.2,
  445.2,
  270.1,
  312.2,
  343.6,
  227.8,
  544.5,
  180.5,
  353.1,
  194.2,
  106.5,
  81.8,
  48.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  18,
  57.2,
  97.9,
  140.5,
  220.7,
  324.2,
  398.6,
  445,
  517.8,
  533.6,
  644.2,
  721,
  717,
  744,
  772,
  811,
  782,
  729,
  715,
  675.2,
  627.8,
  510.6,
  369.2,
  200.3,
  167.3,
  157.5,
  88.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  12.7,
  49.6,
  98,
  155.5,
  224.1,
  298.1,
  374.8,
  448.6,
  519.2,
  588.3,
  655.2,
  669.1,
  689.8,
  745,
  769,
  779,
  776,
  632.3,
  591,
  651,
  592.5,
  509.1,
  412,
  331,
  257.7,
  173.8,
  98,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  13.7,
  59.4,
  121.8,
  194.5,
  267,
  344.8,
  418.4,
  494.7,
  560.9,
  616.5,
  661.8,
  703,
  732,
  744,
  749,
  749,
  731,
  701,
  641.5,
  506.5,
  499.1,
  361.8,
  402.7,
  332.8,
  222.7,
  166.6,
  104.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.1,
  15.2,
  46.1,
  97.4,
  164.2,
  236.5,
  313.5,
  386,
  462.3,
  524.3,
  579.4,
  594.5,
  585.4,
  640.8,
  560.8,
  442.3,
  485,
  436.6,
  470.2,
  500.8,
  385.6,
  429.6,
  348.5,
  241.4,
  155.7,
  151.3,
  122.3,
  67.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  8.1,
  33.5,
  73.6,
  121.1,
  175.8,
  245.8,
  312.5,
  377.3,
  445.7,
  501.4,
  554.2,
  598.9,
  624.5,
  618.6,
  597,
  557.7,
  607.2,
  611.4,
  582.4,
  528.1,
  474.8,
  423.3,
  357.7,
  279.2,
  226.3,
  150.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.2,
  13.5,
  26.9,
  62.4,
  78.7,
  87.6,
  132.3,
  97.6,
  138.8,
  104.3,
  79.7,
  185.8,
  242.3,
  159,
  171.5,
  129.9,
  105.7,
  112.8,
  71.3,
  59.2,
  46.7,
  30.3,
  40,
  38.9,
  22.4,
  24.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.1,
  8.8,
  12.4,
  20.1,
  31.1,
  76.8,
  51.2,
  120.7,
  115.5,
  195.4,
  238.4,
  258.6,
  202.5,
  262.2,
  276.5,
  320.3,
  318.5,
  223.4,
  310.5,
  263.6,
  274.8,
  273.7,
  202.6,
  106,
  55,
  49.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.1,
  32,
  98.5,
  146.3,
  179.6,
  167.4,
  317.3,
  371.8,
  316.8,
  340.6,
  446.7,
  744,
  736,
  677.4,
  677,
  687.3,
  648,
  636.6,
  517.4,
  549.8,
  465.3,
  335.8,
  308.8,
  243.7,
  171.9,
  121.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  8.7,
  44.5,
  50,
  104.1,
  130.6,
  185.3,
  222.4,
  230.5,
  299.2,
  503.4,
  540.3,
  494.7,
  684.8,
  656.4,
  615.1,
  689.2,
  447.9,
  599.2,
  541.7,
  364.1,
  127,
  32.6,
  0,
  2.5,
  3.6,
  65.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.8,
  30.4,
  25.4,
  36.4,
  71.9,
  82.5,
  215.1,
  254.9,
  234.6,
  239,
  215,
  328.2,
  313.2,
  227.5,
  266.3,
  260.6,
  143.7,
  163.5,
  186.7,
  150.6,
  111.9,
  54.2,
  93.7,
  86.9,
  93.4,
  148.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.2,
  19.1,
  40.6,
  59.2,
  86.7,
  97.4,
  181.4,
  200.6,
  289.4,
  402.6,
  433,
  502.8,
  399.4,
  632,
  538.1,
  619.1,
  413.2,
  565.9,
  401,
  365.7,
  107.4,
  94,
  33.8,
  39.7,
  41.6,
  29.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.1,
  16.8,
  9.8,
  30.5,
  47,
  42.6,
  82,
  63.1,
  94.2,
  77.2,
  104.2,
  102.5,
  222.3,
  211.5,
  264.3,
  105.5,
  75.3,
  78,
  118.8,
  194.4,
  131.5,
  125.7,
  177,
  156.7,
  77.7,
  31.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.4,
  20.7,
  56.5,
  134.3,
  183.7,
  177.4,
  219.5,
  210.7,
  272.6,
  247.1,
  322.2,
  256.5,
  439.3,
  209.2,
  171.9,
  378.1,
  335.3,
  348,
  244.6,
  192.2,
  394.3,
  350.8,
  220.2,
  202.1,
  125.1,
  72.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.8,
  19.1,
  46.5,
  63.9,
  117.4,
  126.8,
  191,
  185.2,
  238.1,
  183.4,
  134.2,
  150.1,
  53.2,
  60.8,
  86.8,
  118.7,
  165.4,
  126.9,
  117.5,
  120.2,
  117.2,
  78.8,
  115.5,
  64.5,
  41.4,
  57.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.7,
  12.6,
  30.3,
  82.1,
  170.6,
  184.6,
  387.9,
  454.5,
  578.6,
  592.2,
  585.7,
  659,
  559.8,
  406,
  552.4,
  379.6,
  603.4,
  696.1,
  602.6,
  354,
  181.4,
  269.8,
  186.3,
  224.2,
  204.5,
  117.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.1,
  26.1,
  75.1,
  143.4,
  220.6,
  299,
  351.2,
  361.4,
  470.6,
  507.8,
  427.9,
  538.1,
  541.3,
  562.7,
  658.4,
  602.8,
  469.6,
  574.1,
  629.5,
  471.9,
  342.7,
  114.6,
  119.4,
  82,
  50.2,
  32.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  11.9,
  23.9,
  24.3,
  60,
  121,
  129.6,
  173.4,
  191.6,
  143.2,
  269.3,
  435.5,
  470.2,
  255.7,
  606.6,
  568.8,
  653.6,
  510.7,
  504.9,
  413.5,
  391.7,
  314.1,
  184.3,
  189.6,
  54.5,
  41.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.6,
  23.6,
  63.2,
  137.9,
  188.7,
  277.9,
  346.9,
  425.8,
  492.9,
  552.2,
  612.4,
  525.3,
  552.2,
  732,
  615.2,
  678.4,
  690.9,
  595.7,
  466,
  495.6,
  291.5,
  391.2,
  216.8,
  188.2,
  105.8,
  54.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  9,
  47.2,
  54.4,
  78.4,
  257.6,
  197.9,
  253.6,
  120.3,
  283.6,
  424.9,
  433.4,
  731,
  462.3,
  393.1,
  489.7,
  516.8,
  637.9,
  432.1,
  305.5,
  270.6,
  278.9,
  164.9,
  98.5,
  73.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  15.6,
  40.9,
  57,
  90.3,
  127.6,
  203.2,
  258.3,
  324.5,
  316.4,
  206.3,
  201,
  253.9,
  338.9,
  279.9,
  270,
  386.7,
  321.5,
  391.2,
  308.6,
  237.6,
  89.6,
  131.1,
  80.8,
  46.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  14.5,
  50.3,
  114.7,
  203.1,
  214.9,
  356.2,
  443.5,
  338.2,
  613.4,
  124.5,
  623.8,
  368.8,
  421.1,
  597.2,
  695.7,
  635.5,
  676.5,
  556.6,
  592.6,
  506,
  384.6,
  348.3,
  259.3,
  177.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.6,
  6.9,
  13.1,
  16.3,
  60.9,
  167.9,
  166.4,
  210,
  175.3,
  384.7,
  149.6,
  354.3,
  346.2,
  332.3,
  373.7,
  524.3,
  334.8,
  283.2,
  237.8,
  427.9,
  414.5,
  246.9,
  121.9,
  109.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.3,
  26.3,
  59.4,
  94.7,
  97.9,
  257.1,
  348.4,
  390.6,
  380.6,
  265,
  281.8,
  350,
  402.7,
  389.5,
  388.2,
  492,
  322,
  443,
  276.6,
  262.5,
  160.5,
  66,
  23.6,
  14.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  8.5,
  24.8,
  47,
  84.4,
  128.1,
  194.6,
  280.6,
  296.9,
  333.5,
  353.2,
  414.8,
  445,
  646.5,
  644,
  372.6,
  525.9,
  434.2,
  446.8,
  266.5,
  168.7,
  362.6,
  185.3,
  216.9,
  161.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.9,
  27,
  55.4,
  122.2,
  231.5,
  183.7,
  431.1,
  324.1,
  281.6,
  445.7,
  359.5,
  368.7,
  301.2,
  447,
  414.8,
  590.5,
  592,
  471,
  603.5,
  330.4,
  428.1,
  175.6,
  180.1,
  120.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  11.4,
  39.5,
  85.2,
  118.3,
  191.2,
  303.9,
  451.1,
  461.2,
  323.1,
  435.9,
  477,
  391.1,
  374.5,
  345,
  420.7,
  366.9,
  373.3,
  260.2,
  284.8,
  223.6,
  174.9,
  86.6,
  63.7,
  111.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.4,
  22.8,
  45.2,
  73.8,
  119.5,
  176.9,
  162.3,
  221.6,
  298.9,
  441.6,
  497.4,
  534.3,
  591.3,
  272.4,
  404.7,
  567.7,
  312.2,
  172.1,
  105.7,
  50.4,
  101.4,
  89.9,
  45.7,
  34.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.2,
  56.4,
  119,
  208.6,
  175.5,
  339.4,
  419.3,
  336.9,
  251.2,
  558.4,
  615.3,
  659.3,
  482.1,
  559.2,
  613.9,
  568.3,
  644.4,
  522,
  530.5,
  529.9,
  225.3,
  255.2,
  211.7,
  145.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.4,
  21.5,
  58.6,
  217.7,
  229,
  338.6,
  416.7,
  456.6,
  425.3,
  410.4,
  557.5,
  639,
  691.1,
  364.2,
  493,
  296.4,
  330.1,
  152.8,
  306.3,
  330.2,
  313.9,
  204.2,
  119.1,
  58.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.5,
  38.1,
  88.1,
  165.4,
  239.3,
  350.2,
  365.5,
  435.3,
  400.8,
  445.3,
  465.2,
  610.5,
  547.7,
  474.5,
  484.2,
  441.7,
  420.6,
  431.3,
  322.1,
  306.8,
  279.3,
  213.5,
  171.1,
  113.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3,
  29.5,
  101.9,
  162.9,
  248.3,
  330.1,
  437.8,
  469.8,
  481.7,
  538.7,
  645.4,
  512.8,
  605.1,
  633.8,
  632.2,
  590,
  564.9,
  490.2,
  459.6,
  422.2,
  276.1,
  202.9,
  114.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.4,
  26.4,
  57.2,
  126.1,
  194.6,
  303.9,
  318.6,
  356.9,
  446.8,
  365.4,
  335.1,
  148.5,
  126.7,
  82.5,
  150.7,
  76.9,
  136.2,
  83.1,
  44.8,
  44.5,
  57.3,
  48,
  43.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2,
  17.6,
  49.4,
  96.8,
  168.3,
  228.6,
  251.1,
  241.8,
  283.8,
  404.3,
  355.3,
  224.6,
  446.2,
  563.7,
  547.8,
  532.3,
  441.8,
  362.6,
  245,
  237,
  231.7,
  194.4,
  103,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.7,
  28.2,
  38.1,
  65.8,
  118.7,
  182.6,
  261.8,
  385.6,
  442.2,
  497.8,
  549.1,
  593.5,
  662.1,
  604.7,
  559,
  388.2,
  295.5,
  417.9,
  393.6,
  390.3,
  367.8,
  261.1,
  167,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2,
  37,
  100.8,
  173.6,
  262.5,
  329.1,
  396.2,
  459.4,
  539.5,
  542.5,
  576.1,
  631,
  716,
  519.2,
  344,
  612.6,
  543.3,
  487.7,
  396,
  362.7,
  314.6,
  259.8,
  173,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.6,
  29.9,
  93.9,
  165.2,
  243.1,
  320.1,
  371.8,
  443.3,
  500.9,
  554.9,
  563.8,
  505.9,
  606.7,
  612.8,
  610.7,
  583.1,
  547.6,
  502.7,
  447.8,
  385.5,
  315.6,
  239.9,
  162.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  26.7,
  86,
  157.8,
  236,
  312.4,
  381.8,
  445.3,
  500.9,
  544.9,
  578.3,
  600.5,
  609.4,
  610.6,
  597.3,
  574.7,
  539.6,
  492.9,
  437.9,
  375.4,
  304.5,
  229.4,
  153.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  23.3,
  79.6,
  153.6,
  226.5,
  305.7,
  362.7,
  451.1,
  380.5,
  347.3,
  627.2,
  567.8,
  512.7,
  617.6,
  521.1,
  590.3,
  468.5,
  450,
  296.5,
  178.1,
  76,
  71.8,
  69.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.9,
  16.3,
  34,
  50.7,
  77.2,
  74.4,
  114.3,
  130.6,
  124.9,
  107.4,
  137.9,
  168.3,
  164.4,
  178.6,
  194.4,
  162.7,
  134.4,
  93.9,
  81.2,
  78.2,
  43.6,
  20.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  17.6,
  70.6,
  139.8,
  215.6,
  289.5,
  356.7,
  417.6,
  473.5,
  510.5,
  550.9,
  578.5,
  589.4,
  584.2,
  575,
  544.6,
  504,
  460.9,
  413.9,
  354.5,
  287.9,
  209,
  139.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  13.1,
  54.9,
  119,
  190.6,
  260.8,
  328.4,
  389.7,
  446.1,
  492,
  530.5,
  558.3,
  574.8,
  578.4,
  560.7,
  546.4,
  513.9,
  471.3,
  414.2,
  351.2,
  276.7,
  204.3,
  129.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.5,
  14.4,
  33.6,
  58.6,
  63.2,
  75.5,
  81.3,
  93.1,
  98.9,
  115.1,
  155.8,
  192.2,
  244.3,
  438.7,
  603.8,
  499,
  436.2,
  389.8,
  293.5,
  258.5,
  162.1,
  116.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.1,
  6.7,
  34.6,
  80.8,
  149.3,
  141.8,
  157.8,
  170.1,
  233,
  239.1,
  386.3,
  557.2,
  568.9,
  480.9,
  572.6,
  530.3,
  496.6,
  445.5,
  391,
  328.5,
  255.9,
  178.7,
  103.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.5,
  9.7,
  32.8,
  89.5,
  103.7,
  108.2,
  141.9,
  197.6,
  208.1,
  239.6,
  310.7,
  350.8,
  322,
  406.3,
  291.4,
  237.6,
  303,
  332.8,
  233,
  184.3,
  126.1,
  85.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.7,
  15.4,
  25.5,
  29.4,
  78.4,
  65.4,
  94.5,
  144.2,
  197.4,
  293.9,
  290.7,
  337.9,
  344.3,
  377,
  266.9,
  245.4,
  293.2,
  208.5,
  167.6,
  115.3,
  54.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.4,
  14.5,
  19.7,
  39.8,
  48.3,
  34.9,
  42.5,
  62.1,
  64.6,
  46.8,
  51,
  47.3,
  36.3,
  52.2,
  63.3,
  72.7,
  60.6,
  88.1,
  15.9,
  16.2,
  18.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.6,
  7.2,
  40.2,
  102.1,
  160.7,
  211.2,
  214.2,
  99.9,
  208.4,
  167.8,
  97,
  486.8,
  533.2,
  190.7,
  498.6,
  458.8,
  186.9,
  94,
  105,
  35.1,
  80.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.2,
  16.6,
  41.7,
  66.2,
  193,
  289.7,
  217.1,
  295.2,
  370.1,
  231.7,
  303.7,
  112.4,
  95.5,
  135.2,
  266.9,
  68.5,
  80.2,
  129.2,
  134.8,
  55,
  39,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.5,
  15.2,
  16.4,
  27.8,
  73.3,
  125.5,
  217.3,
  135,
  369.6,
  180.8,
  126.9,
  124.6,
  112.5,
  107.2,
  68.5,
  84.8,
  82.9,
  73.5,
  48.6,
  42.5,
  40.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.1,
  6.5,
  12,
  19.3,
  25.3,
  44.9,
  42.2,
  39.1,
  40.3,
  64.4,
  64.9,
  109.4,
  136.6,
  178.1,
  195.2,
  85.6,
  45.7,
  57.3,
  26.9,
  49.5,
  16.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.9,
  35.3,
  61.8,
  126.7,
  152.6,
  183.7,
  246.3,
  325.1,
  420.7,
  479.4,
  503.8,
  507.8,
  507.9,
  451.5,
  506.2,
  435.8,
  230.8,
  309.5,
  264.4,
  169.6,
  85.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.1,
  2.3,
  14.2,
  19.7,
  17.4,
  35.1,
  49.5,
  66.7,
  114.3,
  214.5,
  249.5,
  404.6,
  266.5,
  317.6,
  36.1,
  195.5,
  272,
  70.8,
  12.6,
  65.8,
  179.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  21.9,
  66.8,
  90.6,
  70.1,
  49,
  37.4,
  40.4,
  48.7,
  33.8,
  60.2,
  45.1,
  64.8,
  52.7,
  87.8,
  81,
  71,
  67.4,
  27.1,
  28.3,
  15.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.4,
  10.3,
  40.5,
  56.2,
  127.1,
  254.9,
  116,
  88.9,
  110.8,
  84.6,
  117,
  98.9,
  102.5,
  103.7,
  99.3,
  49.5,
  65.7,
  50.2,
  37.8,
  27.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.2,
  18.7,
  45.3,
  171.5,
  186.2,
  310.4,
  342.1,
  379.5,
  262.5,
  208,
  294.6,
  176.5,
  148.8,
  204.2,
  460.9,
  213.7,
  197.4,
  247,
  115.1,
  109.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  11.9,
  33.2,
  43.9,
  47.5,
  78.1,
  156.3,
  49,
  190.3,
  524.3,
  277,
  262.4,
  224.1,
  317.7,
  357.3,
  211.4,
  120.1,
  105.1,
  102.6,
  83,
  45.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  11.6,
  41.7,
  135.4,
  251.8,
  244.4,
  328.7,
  303.3,
  215.5,
  212.7,
  161.2,
  185.2,
  400,
  469.5,
  460.8,
  249.4,
  70.2,
  246.4,
  184.2,
  104.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  8.4,
  12.9,
  56.7,
  90.8,
  104.2,
  126.5,
  180.4,
  28.5,
  81.1,
  134.6,
  98.8,
  272.9,
  389.3,
  254.1,
  197.8,
  348.3,
  170.4,
  199.6,
  110.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  13.8,
  53.1,
  100.4,
  52.2,
  209.9,
  269.8,
  308.9,
  254,
  404.4,
  310.5,
  425.3,
  355.5,
  240.9,
  93.1,
  121.3,
  152.6,
  97.4,
  66.9,
  52.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.6,
  8.1,
  30.8,
  50.5,
  78.4,
  76.2,
  65.7,
  99.8,
  94.4,
  150.2,
  173.1,
  186.2,
  155.6,
  212.9,
  169.1,
  152,
  179.9,
  96.4,
  36.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.4,
  6.1,
  24.1,
  46.6,
  67,
  65.7,
  119.5,
  79.9,
  62.2,
  149.4,
  268.3,
  264.6,
  171.2,
  246.8,
  176.2,
  204.3,
  157.6,
  132.9,
  130.7,
  66.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.5,
  7.3,
  15.6,
  24.2,
  42.2,
  133.5,
  124.4,
  117.6,
  154.7,
  176,
  209.7,
  286.5,
  228.7,
  226.4,
  141.5,
  124.2,
  106.9,
  57,
  58.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.5,
  39.4,
  92.3,
  155.6,
  220.1,
  272.9,
  325,
  370,
  404.7,
  426,
  435.7,
  435.7,
  423.2,
  397.6,
  358.7,
  314.9,
  262,
  206.9,
  142.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.9,
  38,
  114.7,
  122.3,
  137.6,
  227.2,
  303.6,
  330.4,
  386.7,
  407.6,
  404.3,
  423,
  418.1,
  388.2,
  353.8,
  303.9,
  242.5,
  183.6,
  116.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  4,
  12.2,
  29.2,
  43,
  58.4,
  77.1,
  124.2,
  157.1,
  174.9,
  106.7,
  142.5,
  162.7,
  219.8,
  293.3,
  385,
  352.3,
  159.4,
  120.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.2,
  28.6,
  31.1,
  146.7,
  228.7,
  307.2,
  358.4,
  228.8,
  234.5,
  446.1,
  452.4,
  452,
  436.4,
  411,
  379.1,
  330.7,
  248.1,
  189,
  120.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.5,
  32.7,
  90.2,
  155.7,
  221.4,
  281,
  333.9,
  374.9,
  409.3,
  431.2,
  443.6,
  449.1,
  438.5,
  411.7,
  376.4,
  325.4,
  269.3,
  208.8,
  140.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.8,
  12.6,
  28.4,
  44,
  63,
  73.1,
  85.3,
  94.4,
  158.2,
  258.3,
  356.6,
  57.7,
  160.3,
  170.2,
  197.3,
  135.9,
  69.4,
  135.9,
  40.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.7,
  24.8,
  87.4,
  171.8,
  138.3,
  153.7,
  156.7,
  230.1,
  377.8,
  293.7,
  173.4,
  446,
  195.1,
  283.8,
  314.3,
  168.4,
  146.3,
  165.5,
  98.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.7,
  10.8,
  24.5,
  38.6,
  54,
  52.2,
  62.9,
  147.9,
  101.5,
  29.3,
  116.9,
  150.3,
  279.6,
  89.2,
  45.2,
  28.7,
  85.5,
  50,
  11,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.1,
  12.6,
  36.3,
  78.4,
  136.5,
  166.2,
  291.2,
  326,
  279.1,
  358.9,
  283.3,
  271.5,
  199,
  158,
  63,
  84.2,
  49.3,
  37.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  23.9,
  78.8,
  144.5,
  205,
  271.4,
  325.7,
  368.4,
  401.9,
  425.4,
  434.8,
  432.5,
  414.5,
  386.9,
  348.8,
  301,
  243.1,
  178.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  20.9,
  76.5,
  141.4,
  205.6,
  264.8,
  315.8,
  358.9,
  391.7,
  413.2,
  424.1,
  423.2,
  404.6,
  378.5,
  339.7,
  292,
  234.1,
  169,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  25.3,
  79.7,
  133.4,
  191.5,
  226.4,
  254.1,
  331.8,
  389.3,
  398.6,
  387.4,
  432.3,
  371.5,
  257.1,
  277.7,
  232.4,
  148.1,
  108.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  11.8,
  29.7,
  53.5,
  83.4,
  117.9,
  148.5,
  166.7,
  186.4,
  224.4,
  307.8,
  316.4,
  285.3,
  221.3,
  171,
  128.4,
  105.4,
  78.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  13.9,
  58.9,
  117.8,
  179.7,
  238.4,
  290.2,
  332.5,
  362.8,
  381.6,
  388.6,
  387.1,
  369.7,
  345,
  310.5,
  263.5,
  210.1,
  149.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.2,
  13.8,
  23.4,
  34.6,
  57.5,
  59.3,
  73.4,
  92.6,
  100.4,
  105.1,
  119.3,
  151.5,
  192,
  216,
  211.2,
  172.6,
  72.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.1,
  6.2,
  20.2,
  34.6,
  63.7,
  93,
  111.2,
  134.6,
  176.1,
  108.9,
  82,
  79.8,
  76.2,
  90.3,
  89.7,
  61,
  33.3,
  23.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.1,
  8.7,
  19.5,
  38.9,
  66.8,
  71.8,
  79.8,
  130.9,
  158.1,
  197.6,
  159.8,
  83,
  45.5,
  31.1,
  29.4,
  46.7,
  43.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.3,
  42.9,
  98.2,
  154.1,
  212,
  262.4,
  303.9,
  335.6,
  353.9,
  363,
  360.5,
  344,
  319,
  282.5,
  236.6,
  186.4,
  112.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.7,
  12.2,
  22.1,
  98.8,
  155.1,
  76.9,
  112.7,
  172.6,
  233.7,
  310.2,
  334.5,
  219.7,
  128.2,
  116.6,
  145.2,
  43.9,
  23.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.1,
  8.3,
  9.7,
  49.3,
  46.3,
  108.5,
  135.4,
  122.9,
  127.5,
  119.6,
  106.8,
  90.1,
  162.5,
  111,
  79.7,
  28.6,
  57.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.7,
  15,
  17.5,
  21.6,
  19.2,
  27.2,
  37.2,
  31.1,
  19.1,
  16,
  14.8,
  11.8,
  10.8,
  9.6,
  9.8,
  5.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.1,
  20.5,
  64.5,
  68.4,
  47.2,
  53,
  69,
  187.4,
  108.4,
  80.9,
  207.6,
  87.8,
  57.1,
  115.6,
  163.5,
  145.7,
  76.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.4,
  8.2,
  42,
  128.3,
  185.3,
  225.4,
  258.1,
  270.4,
  315.3,
  312.8,
  237,
  247.8,
  167.8,
  119.8,
  153.7,
  163.7,
  95.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.7,
  7.5,
  26,
  24.8,
  21.4,
  29.4,
  40.9,
  88.1,
  158.3,
  79.2,
  207.4,
  143.5,
  220.9,
  214.5,
  133.3,
  66.3,
  31.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.2,
  20.8,
  26,
  32.1,
  44.7,
  69.1,
  85.5,
  38,
  73.8,
  68.1,
  52.3,
  40,
  25.1,
  48,
  48.3,
  33.2,
  9.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.9,
  27.6,
  67.7,
  97.1,
  111,
  112.8,
  208.8,
  163.3,
  132.8,
  124.2,
  151.9,
  155.1,
  121.9,
  92.9,
  60.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.6,
  9.3,
  19.8,
  39.4,
  64.6,
  70.2,
  74.3,
  87.5,
  105.3,
  104.8,
  93.8,
  79.8,
  66.7,
  68.6,
  48.5,
  35.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  14.6,
  34,
  92.4,
  136.7,
  149,
  240.8,
  121.9,
  176.2,
  108.6,
  64.3,
  53.1,
  40.9,
  30,
  20.9,
  15.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.7,
  3.8,
  6.8,
  10.4,
  19.4,
  21.7,
  28.5,
  25.8,
  29.5,
  28.2,
  21.3,
  23.9,
  35.7,
  18.9,
  10.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.4,
  9.9,
  25.6,
  40.6,
  55.5,
  74.5,
  72,
  59.4,
  59.6,
  59.5,
  46,
  36.2,
  33.4,
  39.1,
  39.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.6,
  11.1,
  50.7,
  101.7,
  153.3,
  200.6,
  241.5,
  268.6,
  292,
  294.8,
  296.6,
  264,
  182.6,
  154.8,
  107.2,
  81.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  9.8,
  46,
  95.3,
  149.4,
  200.6,
  242.4,
  259.3,
  263.7,
  276.5,
  301.9,
  276.6,
  260.6,
  224.5,
  178.5,
  109.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  9.3,
  39.3,
  84.3,
  133.6,
  182.5,
  221.6,
  253,
  276.7,
  289.8,
  291.5,
  279.5,
  255.9,
  219.9,
  177.2,
  126.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.1,
  4.8,
  13.7,
  25.9,
  39.7,
  30.4,
  77.7,
  76.5,
  100.4,
  135.2,
  208.2,
  69.8,
  43.2,
  63.4,
  20.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.3,
  18.9,
  56.9,
  78.9,
  72.9,
  76.7,
  90.1,
  98.9,
  38.2,
  82.7,
  89,
  44.5,
  18.6,
  16.7,
  16.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.1,
  12.4,
  28.5,
  53.5,
  61.3,
  58.3,
  101.3,
  101.3,
  81.6,
  65.5,
  40.9,
  41.8,
  88.5,
  55.3,
  45,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.8,
  8,
  10.7,
  12.5,
  29.6,
  58.8,
  46.4,
  53.2,
  58,
  74.4,
  67.9,
  41.4,
  25.2,
  19.6,
  30.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.5,
  7.5,
  17.6,
  24.1,
  49.3,
  60.4,
  55.9,
  59.6,
  74.9,
  125.2,
  97.6,
  101,
  84.7,
  62.1,
  32.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.7,
  21,
  28.9,
  49.9,
  99.2,
  207.3,
  183.5,
  146.3,
  146.7,
  158.7,
  163.5,
  199.5,
  163,
  140.8,
  95.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.8,
  18,
  38,
  48.1,
  61.5,
  69.4,
  79.2,
  92.8,
  117.8,
  123.4,
  93.3,
  146.6,
  96.2,
  64.9,
  29.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.5,
  4,
  8,
  15.3,
  26,
  37.7,
  56.8,
  59.6,
  52.7,
  57.2,
  33.9,
  32.7,
  27.1,
  18.4,
  13.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.7,
  3.9,
  14.7,
  13.4,
  17.9,
  37.5,
  48.1,
  48.6,
  59.2,
  81.4,
  55,
  29.6,
  26.4,
  27.8,
  26.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  10.9,
  20.1,
  27.5,
  46.2,
  73.2,
  31.9,
  59.2,
  82.9,
  48.1,
  68.4,
  70.7,
  76.7,
  35.4,
  26.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.2,
  7.1,
  11.9,
  25.3,
  50.4,
  45.7,
  46.1,
  29.4,
  30.1,
  21.1,
  14.4,
  11,
  12.9,
  10.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.1,
  17.9,
  69.1,
  176,
  178.1,
  171.8,
  214.5,
  239.2,
  250.3,
  249.2,
  225.9,
  72.6,
  194.4,
  110.5,
  43.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  9.8,
  19.4,
  33.1,
  48,
  67.1,
  79.7,
  73.2,
  76.8,
  74.8,
  84,
  90.4,
  67.9,
  46.3,
  31.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  8.4,
  24.8,
  49,
  74.4,
  97.3,
  142.4,
  204.9,
  235.5,
  246.4,
  213.5,
  171.3,
  77.6,
  62,
  40.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.7,
  39.6,
  63.4,
  109.7,
  84.9,
  64.5,
  56.1,
  33,
  19.8,
  16,
  25.9,
  16.7,
  13.1,
  11.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.6,
  6,
  20.4,
  29.8,
  19.5,
  20.1,
  48.5,
  87.6,
  52.5,
  93.5,
  206.2,
  187.5,
  157.8,
  91.6,
  33.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.4,
  19.9,
  23.9,
  28.8,
  45.5,
  36,
  23,
  28.1,
  22.2,
  16.6,
  12.5,
  8.3,
  7.3,
  4.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.9,
  24.1,
  46,
  37.5,
  33,
  39.4,
  47.1,
  49.3,
  42.8,
  53.3,
  40.7,
  74.7,
  77,
  53.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.9,
  6,
  11.5,
  18.5,
  29.4,
  44,
  46.8,
  45.4,
  47,
  51.3,
  37.2,
  22.8,
  18.1,
  9.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  6.1,
  12.2,
  27.1,
  33.4,
  82.8,
  82,
  94.5,
  173.2,
  164.1,
  91.8,
  72,
  64.1,
  39.2,
  74.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.1,
  8.9,
  22.2,
  17.9,
  18.6,
  16.7,
  17.8,
  16.8,
  18.5,
  17,
  10.8,
  5.8,
  9.9,
  9.9,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.8,
  6.7,
  7.4,
  7.4,
  10.6,
  16.1,
  11.5,
  74.1,
  56.3,
  67.6,
  96.3,
  68.2,
  59.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.5,
  9.1,
  14.1,
  53.7,
  62.5,
  76,
  89.8,
  60,
  69.1,
  42.2,
  18.1,
  27.7,
  37.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  7.7,
  24.3,
  67.7,
  81.7,
  141.2,
  182.8,
  200.7,
  225.3,
  194.8,
  142.6,
  89.3,
  58,
  25,
  20.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.2,
  31.1,
  40.4,
  44.6,
  136,
  192.5,
  217.8,
  149.1,
  130.6,
  209.1,
  105.1,
  96.9,
  49,
  70.5,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  3.5,
  7.7,
  11.2,
  15.7,
  37.6,
  33.9,
  42.7,
  68.2,
  78.7,
  83.5,
  74,
  66.2,
  88,
  46.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.9,
  19.5,
  32.7,
  66.9,
  120.7,
  128,
  147.6,
  114.7,
  189.3,
  200,
  179.9,
  154.2,
  115.2,
  74.3,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  4.1,
  24.9,
  41.4,
  108.5,
  141.6,
  173.9,
  181.7,
  182.5,
  59.5,
  104.6,
  68.3,
  38.4,
  35,
  26.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  5.8,
  32.2,
  56.2,
  67.5,
  67.2,
  69,
  65.8,
  66.6,
  38.5,
  13.2,
  27,
  38.2,
  22.6,
  9.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.1,
  5.6,
  17.5,
  38.3,
  80.2,
  53.2,
  28.9,
  85.8,
  101.8,
  118.2,
  129.7,
  38.7,
  50.6,
  21.6,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.1,
  11.8,
  25,
  50,
  82.2,
  92.2,
  112.9,
  124.6,
  123.6,
  124.5,
  124.7,
  119.2,
  120.9,
  61.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  3.5,
  14.9,
  23.7,
  26.3,
  31.2,
  31.2,
  24.3,
  26.5,
  25.3,
  27,
  25.2,
  16.9,
  12.2,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.9,
  5.6,
  10.7,
  18.7,
  36,
  44.5,
  37,
  38.5,
  28.9,
  29.6,
  26.6,
  20.5,
  17.7,
  11.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.6,
  5.8,
  15,
  21.2,
  23.8,
  32.8,
  32.9,
  33.2,
  31.4,
  34.2,
  43.1,
  49.8,
  25.3,
  17.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.3,
  2.5,
  7.4,
  10,
  16.8,
  16.7,
  17,
  14.1,
  13,
  10.8,
  9.1,
  9.2,
  7.8,
  6.1,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.6,
  9.6,
  34.3,
  57.6,
  100.9,
  102.2,
  90.9,
  76,
  39,
  21.1,
  14,
  14.3,
  12.9,
  5.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  10.8,
  21.6,
  12.4,
  13.2,
  16.2,
  44.2,
  39.2,
  67,
  49.4,
  13.3,
  15.4,
  7.3,
  12.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.8,
  12.6,
  36,
  53,
  56.1,
  57.4,
  46.9,
  32.6,
  52.2,
  42.6,
  36,
  21.6,
  69.4,
  16.7,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.3,
  21.8,
  76.9,
  96.5,
  111.2,
  86.1,
  143.5,
  154.1,
  164.9,
  158.2,
  83.1,
  106.8,
  114.5,
  40.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.8,
  19.9,
  50.6,
  111.3,
  132.2,
  162.5,
  198.4,
  216.6,
  215.3,
  209.1,
  153.3,
  83.9,
  72,
  46.4,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  1.2,
  14.3,
  31.5,
  66.2,
  145.6,
  128.1,
  158.4,
  91,
  95.2,
  91.3,
  86.4,
  100.1,
  118.2,
  39,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  2.2,
  5.4,
  10,
  16,
  17.4,
  24.3,
  27.7,
  20.1,
  16.5,
  29.4,
  50.6,
  49.2,
  32.8,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 Tair =
  259.8,     259.8,   259.8,   259.8, 
  259.7,     259.7,   259.7,   259.7,
  259.6,     259.6,   259.6,   259.6,
  259.5,     259.5,   259.5,   259.5,
  259.4,     259.4,   259.4,   259.4,
  259.35,    259.35,  259.35,  259.35,
  259.3,     259.3,   259.3,   259.3,
  259.25,    259.25,  259.25,  259.25,
  259.15,    259.15,  259.15,  259.15,
  258.95,    258.95,  258.95,  258.95,
  258.8,     258.8,   258.8,   258.8,
  258.75,    258.75,  258.75,  258.75,
  258.75,    258.75,  258.75,  258.75,
  258.85,    258.85,  258.85,  258.85,
  258.9,     258.9,   258.9,   258.9,
  258.9,     258.9,   258.9,   258.9,
  259,       259,     259,     259,
  259.1,     259.1,   259.1,   259.1,
  259.2,     259.2,   259.2,   259.2,
  259.45,    259.45,  259.45,  259.45,
  259.85,    259.85,  259.85,  259.85,
  260.3,     260.3,   260.3,   260.3,
  260.85,    260.85,  260.85,  260.85,
  261.45,    261.45,  261.45,  261.45,
  262.1,     262.1,   262.1,   262.1,
  262.65,    262.65,  262.65,  262.65,
  263.1,     263.1,   263.1,   263.1,
  263.45,    263.45,  263.45,  263.45,
  263.6,     263.6,   263.6,   263.6,
  263.55,    263.55,  263.55,  263.55,
  263.45,    263.45,  263.45,  263.45,
  263.4,     263.4,   263.4,   263.4,
  263.1,     263.1,   263.1,   263.1,
  262.5,     262.5,   262.5,   262.5,
  261.85,    261.85,  261.85,  261.85,
  261.25,    261.25,  261.25,  261.25,
  260.9,     260.9,   260.9,   260.9,
  260.85,    260.85,  260.85,  260.85,
  260.75,    260.75,  260.75,  260.75,
  260.5,     260.5,   260.5,   260.5,
  260.2,     260.2,   260.2,   260.2,
  259.85,    259.85,  259.85,  259.85,
  259.35,    259.35,  259.35,  259.35,
  258.9,     258.9,   258.9,   258.9,
  258.7,     258.7,   258.7,   258.7,
  258.5,     258.5,   258.5,   258.5,
  258.2,     258.2,   258.2,   258.2,
  258.05,    258.05,  258.05,  258.05,
  257.8,     257.8,   257.8,   257.8,
  257.5,     257.5,   257.5,   257.5,
  257.4,     257.4,   257.4,   257.4,
  257.35,    257.35,  257.35,  257.35,
  257.3,     257.3,   257.3,   257.3,
  257.2,     257.2,   257.2,   257.2,
  257,       257,     257,     257,
  256.75,    256.75,  256.75,  256.75,
  256.5,     256.5,   256.5,   256.5,
  256.4,     256.4,   256.4,   256.4,
  256.25,    256.25,  256.25,  256.25,
  255.95,    255.95,  255.95,  255.95,
  255.9,     255.9,   255.9,   255.9,
  255.9,     255.9,   255.9,   255.9,
  255.85,    255.85,  255.85,  255.85,
  255.85,    255.85,  255.85,  255.85,
  255.8,     255.8,   255.8,   255.8,
  255.8,     255.8,   255.8,   255.8,
  255.85,    255.85,  255.85,  255.85,
  256.25,    256.25,  256.25,  256.25,
  257,       257,     257,     257,
  258,       258,     258,     258,
  259.2,     259.2,   259.2,   259.2,
  260.15,    260.15,  260.15,  260.15,
  260.95,    260.95,  260.95,  260.95,
  261.8,     261.8,   261.8,   261.8,
  262.65,    262.65,  262.65,  262.65,
  263.2,     263.2,   263.2,   263.2,
  263.5,     263.5,   263.5,   263.5,
  263.6,     263.6,   263.6,   263.6,
  263.55,    263.55,  263.55,  263.55,
  263.35,    263.35,  263.35,  263.35,
  262.85,    262.85,  262.85,  262.85,
  262.2,     262.2,   262.2,   262.2,
  261.6,     261.6,   261.6,   261.6,
  261.15,    261.15,  261.15,  261.15,
  260.75,    260.75,  260.75,  260.75,
  260.45,    260.45,  260.45,  260.45,
  260.3,     260.3,   260.3,   260.3,
  260.2,     260.2,   260.2,   260.2,
  260.1,     260.1,   260.1,   260.1,
  260.05,    260.05,  260.05,  260.05,
  260.05,    260.05,  260.05,  260.05,
  260.05,    260.05,  260.05,  260.05,
  260,       260,     260,     260,
  259.9,     259.9,   259.9,   259.9,
  259.85,    259.85,  259.85,  259.85,
  259.9,     259.9,   259.9,   259.9,
  260.05,    260.05,  260.05,  260.05,
  260.2,     260.2,   260.2,   260.2,
  260.45,    260.45,  260.45,  260.45,
  260.9,     260.9,   260.9,   260.9,
  261.25,    261.25,  261.25,  261.25,
  261.25,    261.25,  261.25,  261.25,
  261.15,    261.15,  261.15,  261.15,
  261.1,     261.1,   261.1,   261.1,
  261.1,     261.1,   261.1,   261.1,
  261.3,     261.3,   261.3,   261.3,
  261.5,     261.5,   261.5,   261.5,
  261.6,     261.6,   261.6,   261.6,
  261.8,     261.8,   261.8,   261.8,
  262.1,     262.1,   262.1,   262.1,
  262.25,    262.25,  262.25,  262.25,
  262.35,    262.35,  262.35,  262.35,
  262.6,     262.6,   262.6,   262.6,
  262.9,     262.9,   262.9,   262.9,
  263.25,    263.25,  263.25,  263.25,
  263.55,    263.55,  263.55,  263.55,
  263.8,     263.8,   263.8,   263.8,
  264.15,    264.15,  264.15,  264.15,
  264.55,    264.55,  264.55,  264.55,
  265,       265,     265,     265,
  265.45,    265.45,  265.45,  265.45,
  265.75,    265.75,  265.75,  265.75,
  265.95,    265.95,  265.95,  265.95,
  266.15,    266.15,  266.15,  266.15,
  266.35,    266.35,  266.35,  266.35,
  266.55,    266.55,  266.55,  266.55,
  266.6,     266.6,   266.6,   266.6,
  266.6,     266.6,   266.6,   266.6,
  266.7,     266.7,   266.7,   266.7,
  266.75,    266.75,  266.75,  266.75,
  266.7,     266.7,   266.7,   266.7,
  266.65,    266.65,  266.65,  266.65,
  266.55,    266.55,  266.55,  266.55,
  266.5,     266.5,   266.5,   266.5,
  266.6,     266.6,   266.6,   266.6,
  266.75,    266.75,  266.75,  266.75,
  266.85,    266.85,  266.85,  266.85,
  266.85,    266.85,  266.85,  266.85,
  266.85,    266.85,  266.85,  266.85,
  266.9,     266.9,   266.9,   266.9,
  267.05,    267.05,  267.05,  267.05,
  267.25,    267.25,  267.25,  267.25,
  267.4,     267.4,   267.4,   267.4,
  267.45,    267.45,  267.45,  267.45,
  267.5,     267.5,   267.5,   267.5,
  267.55,    267.55,  267.55,  267.55,
  267.55,    267.55,  267.55,  267.55,
  267.55,    267.55,  267.55,  267.55,
  267.6,     267.6,   267.6,   267.6,
  267.7,     267.7,   267.7,   267.7,
  267.75,    267.75,  267.75,  267.75,
  267.75,    267.75,  267.75,  267.75,
  267.75,    267.75,  267.75,  267.75,
  267.75,    267.75,  267.75,  267.75,
  267.75,    267.75,  267.75,  267.75,
  267.75,    267.75,  267.75,  267.75,
  267.75,    267.75,  267.75,  267.75,
  267.65,    267.65,  267.65,  267.65,
  267.55,    267.55,  267.55,  267.55,
  267.5,     267.5,   267.5,   267.5,
  267.4,     267.4,   267.4,   267.4,
  267.4,     267.4,   267.4,   267.4,
  267.4,     267.4,   267.4,   267.4,
  267.3,     267.3,   267.3,   267.3,
  267.2,     267.2,   267.2,   267.2,
  267.2,     267.2,   267.2,   267.2,
  267.3,     267.3,   267.3,   267.3,
  267.35,    267.35,  267.35,  267.35,
  267.45,    267.45,  267.45,  267.45,
  267.65,    267.65,  267.65,  267.65,
  267.85,    267.85,  267.85,  267.85,
  268,       268,     268,     268,
  268.15,    268.15,  268.15,  268.15,
  268.25,    268.25,  268.25,  268.25,
  268.3,     268.3,   268.3,   268.3,
  268.35,    268.35,  268.35,  268.35,
  268.35,    268.35,  268.35,  268.35,
  268.4,     268.4,   268.4,   268.4,
  268.45,    268.45,  268.45,  268.45,
  268.5,     268.5,   268.5,   268.5,
  268.65,    268.65,  268.65,  268.65,
  268.85,    268.85,  268.85,  268.85,
  269.05,    269.05,  269.05,  269.05,
  269.2,     269.2,   269.2,   269.2,
  269.3,     269.3,   269.3,   269.3,
  269.35,    269.35,  269.35,  269.35,
  269.35,    269.35,  269.35,  269.35,
  269.2,     269.2,   269.2,   269.2,
  268.95,    268.95,  268.95,  268.95,
  268.85,    268.85,  268.85,  268.85,
  268.85,    268.85,  268.85,  268.85,
  268.8,     268.8,   268.8,   268.8,
  268.7,     268.7,   268.7,   268.7,
  268.5,     268.5,   268.5,   268.5,
  268.4,     268.4,   268.4,   268.4,
  268.5,     268.5,   268.5,   268.5,
  268.55,    268.55,  268.55,  268.55,
  268.45,    268.45,  268.45,  268.45,
  268.3,     268.3,   268.3,   268.3,
  268.25,    268.25,  268.25,  268.25,
  268.15,    268.15,  268.15,  268.15,
  267.9,     267.9,   267.9,   267.9,
  267.55,    267.55,  267.55,  267.55,
  267.2,     267.2,   267.2,   267.2,
  267.15,    267.15,  267.15,  267.15,
  267.2,     267.2,   267.2,   267.2,
  267.25,    267.25,  267.25,  267.25,
  267.4,     267.4,   267.4,   267.4,
  267.5,     267.5,   267.5,   267.5,
  267.55,    267.55,  267.55,  267.55,
  267.55,    267.55,  267.55,  267.55,
  267.6,     267.6,   267.6,   267.6,
  267.75,    267.75,  267.75,  267.75,
  268.05,    268.05,  268.05,  268.05,
  268.45,    268.45,  268.45,  268.45,
  268.7,     268.7,   268.7,   268.7,
  268.65,    268.65,  268.65,  268.65,
  268.4,     268.4,   268.4,   268.4,
  268.4,     268.4,   268.4,   268.4,
  268.7,     268.7,   268.7,   268.7,
  268.75,    268.75,  268.75,  268.75,
  268.8,     268.8,   268.8,   268.8,
  269.05,    269.05,  269.05,  269.05,
  269.15,    269.15,  269.15,  269.15,
  269,       269,     269,     269,
  268.45,    268.45,  268.45,  268.45,
  267.65,    267.65,  267.65,  267.65,
  267.05,    267.05,  267.05,  267.05,
  266.65,    266.65,  266.65,  266.65,
  266.15,    266.15,  266.15,  266.15,
  265.55,    265.55,  265.55,  265.55,
  265,       265,     265,     265,
  264.5,     264.5,   264.5,   264.5,
  264.2,     264.2,   264.2,   264.2,
  264.15,    264.15,  264.15,  264.15,
  263.95,    263.95,  263.95,  263.95,
  263.6,     263.6,   263.6,   263.6,
  263.25,    263.25,  263.25,  263.25,
  263.25,    263.25,  263.25,  263.25,
  263.55,    263.55,  263.55,  263.55,
  263.7,     263.7,   263.7,   263.7,
  263.6,     263.6,   263.6,   263.6,
  263.35,    263.35,  263.35,  263.35,
  263.5,     263.5,   263.5,   263.5,
  264.05,    264.05,  264.05,  264.05,
  264.65,    264.65,  264.65,  264.65,
  265.4,     265.4,   265.4,   265.4,
  266.15,    266.15,  266.15,  266.15,
  266.55,    266.55,  266.55,  266.55,
  266.65,    266.65,  266.65,  266.65,
  266.55,    266.55,  266.55,  266.55,
  266.45,    266.45,  266.45,  266.45,
  266.35,    266.35,  266.35,  266.35,
  266.15,    266.15,  266.15,  266.15,
  266,       266,     266,     266,
  265.9,     265.9,   265.9,   265.9,
  265.85,    265.85,  265.85,  265.85,
  265.9,     265.9,   265.9,   265.9,
  265.85,    265.85,  265.85,  265.85,
  265.5,     265.5,   265.5,   265.5,
  265.2,     265.2,   265.2,   265.2,
  265.05,    265.05,  265.05,  265.05,
  264.9,     264.9,   264.9,   264.9,
  264.95,    264.95,  264.95,  264.95,
  265.15,    265.15,  265.15,  265.15,
  265.15,    265.15,  265.15,  265.15,
  265.15,    265.15,  265.15,  265.15,
  265.3,     265.3,   265.3,   265.3,
  265.35,    265.35,  265.35,  265.35,
  265.4,     265.4,   265.4,   265.4,
  265.35,    265.35,  265.35,  265.35,
  265.15,    265.15,  265.15,  265.15,
  264.95,    264.95,  264.95,  264.95,
  264.7,     264.7,   264.7,   264.7,
  264.4,     264.4,   264.4,   264.4,
  264.25,    264.25,  264.25,  264.25,
  264.25,    264.25,  264.25,  264.25,
  264.25,    264.25,  264.25,  264.25,
  264.2,     264.2,   264.2,   264.2,
  264.05,    264.05,  264.05,  264.05,
  263.9,     263.9,   263.9,   263.9,
  263.95,    263.95,  263.95,  263.95,
  264.35,    264.35,  264.35,  264.35,
  264.9,     264.9,   264.9,   264.9,
  265.35,    265.35,  265.35,  265.35,
  265.75,    265.75,  265.75,  265.75,
  266,       266,     266,     266,
  266.15,    266.15,  266.15,  266.15,
  266.3,     266.3,   266.3,   266.3,
  266.4,     266.4,   266.4,   266.4,
  266.45,    266.45,  266.45,  266.45,
  266.5,     266.5,   266.5,   266.5,
  266.6,     266.6,   266.6,   266.6,
  266.75,    266.75,  266.75,  266.75,
  266.95,    266.95,  266.95,  266.95,
  267.15,    267.15,  267.15,  267.15,
  267.3,     267.3,   267.3,   267.3,
  267.45,    267.45,  267.45,  267.45,
  267.6,     267.6,   267.6,   267.6,
  267.7,     267.7,   267.7,   267.7,
  267.8,     267.8,   267.8,   267.8,
  267.9,     267.9,   267.9,   267.9,
  268.05,    268.05,  268.05,  268.05,
  268.2,     268.2,   268.2,   268.2,
  268.2,     268.2,   268.2,   268.2,
  268.05,    268.05,  268.05,  268.05,
  267.95,    267.95,  267.95,  267.95,
  268,       268,     268,     268,
  268.1,     268.1,   268.1,   268.1,
  268.25,    268.25,  268.25,  268.25,
  268.4,     268.4,   268.4,   268.4,
  268.5,     268.5,   268.5,   268.5,
  268.55,    268.55,  268.55,  268.55,
  268.55,    268.55,  268.55,  268.55,
  268.55,    268.55,  268.55,  268.55,
  268.65,    268.65,  268.65,  268.65,
  268.85,    268.85,  268.85,  268.85,
  269,       269,     269,     269,
  269,       269,     269,     269,
  268.95,    268.95,  268.95,  268.95,
  268.8,     268.8,   268.8,   268.8,
  268.45,    268.45,  268.45,  268.45,
  268.1,     268.1,   268.1,   268.1,
  267.8,     267.8,   267.8,   267.8,
  267.5,     267.5,   267.5,   267.5,
  267.05,    267.05,  267.05,  267.05,
  266.35,    266.35,  266.35,  266.35,
  265.85,    265.85,  265.85,  265.85,
  265.65,    265.65,  265.65,  265.65,
  265.35,    265.35,  265.35,  265.35,
  265.35,    265.35,  265.35,  265.35,
  265.8,     265.8,   265.8,   265.8,
  266.2,     266.2,   266.2,   266.2,
  266.3,     266.3,   266.3,   266.3,
  266.15,    266.15,  266.15,  266.15,
  266.05,    266.05,  266.05,  266.05,
  266.05,    266.05,  266.05,  266.05,
  266.05,    266.05,  266.05,  266.05,
  266,       266,     266,     266,
  265.8,     265.8,   265.8,   265.8,
  265.55,    265.55,  265.55,  265.55,
  265.4,     265.4,   265.4,   265.4,
  265.25,    265.25,  265.25,  265.25,
  265.05,    265.05,  265.05,  265.05,
  264.9,     264.9,   264.9,   264.9,
  264.8,     264.8,   264.8,   264.8,
  264.75,    264.75,  264.75,  264.75,
  264.7,     264.7,   264.7,   264.7,
  264.55,    264.55,  264.55,  264.55,
  264.4,     264.4,   264.4,   264.4,
  264.3,     264.3,   264.3,   264.3,
  264.3,     264.3,   264.3,   264.3,
  264.4,     264.4,   264.4,   264.4,
  264.5,     264.5,   264.5,   264.5,
  264.6,     264.6,   264.6,   264.6,
  264.65,    264.65,  264.65,  264.65,
  264.7,     264.7,   264.7,   264.7,
  264.8,     264.8,   264.8,   264.8,
  264.85,    264.85,  264.85,  264.85,
  264.85,    264.85,  264.85,  264.85,
  264.9,     264.9,   264.9,   264.9,
  265.05,    265.05,  265.05,  265.05,
  265.25,    265.25,  265.25,  265.25,
  265.4,     265.4,   265.4,   265.4,
  265.45,    265.45,  265.45,  265.45,
  265.55,    265.55,  265.55,  265.55,
  265.7,     265.7,   265.7,   265.7,
  265.75,    265.75,  265.75,  265.75,
  265.6,     265.6,   265.6,   265.6,
  265.4,     265.4,   265.4,   265.4,
  265.1,     265.1,   265.1,   265.1,
  264.8,     264.8,   264.8,   264.8,
  264.8,     264.8,   264.8,   264.8,
  264.75,    264.75,  264.75,  264.75,
  264.6,     264.6,   264.6,   264.6,
  264.5,     264.5,   264.5,   264.5,
  264.35,    264.35,  264.35,  264.35,
  264.2,     264.2,   264.2,   264.2,
  264.2,     264.2,   264.2,   264.2,
  264.25,    264.25,  264.25,  264.25,
  264.25,    264.25,  264.25,  264.25,
  264.15,    264.15,  264.15,  264.15,
  264,       264,     264,     264,
  263.85,    263.85,  263.85,  263.85,
  263.75,    263.75,  263.75,  263.75,
  263.7,     263.7,   263.7,   263.7,
  263.65,    263.65,  263.65,  263.65,
  263.6,     263.6,   263.6,   263.6,
  263.55,    263.55,  263.55,  263.55,
  263.6,     263.6,   263.6,   263.6,
  263.6,     263.6,   263.6,   263.6,
  263.55,    263.55,  263.55,  263.55,
  263.55,    263.55,  263.55,  263.55,
  263.5,     263.5,   263.5,   263.5,
  263.45,    263.45,  263.45,  263.45,
  263.4,     263.4,   263.4,   263.4,
  263.3,     263.3,   263.3,   263.3,
  263.2,     263.2,   263.2,   263.2,
  263.25,    263.25,  263.25,  263.25,
  263.55,    263.55,  263.55,  263.55,
  263.95,    263.95,  263.95,  263.95,
  264.25,    264.25,  264.25,  264.25,
  264.4,     264.4,   264.4,   264.4,
  264.45,    264.45,  264.45,  264.45,
  264.5,     264.5,   264.5,   264.5,
  264.65,    264.65,  264.65,  264.65,
  264.85,    264.85,  264.85,  264.85,
  265.1,     265.1,   265.1,   265.1,
  265.35,    265.35,  265.35,  265.35,
  265.6,     265.6,   265.6,   265.6,
  265.8,     265.8,   265.8,   265.8,
  265.85,    265.85,  265.85,  265.85,
  265.95,    265.95,  265.95,  265.95,
  266.05,    266.05,  266.05,  266.05,
  266.05,    266.05,  266.05,  266.05,
  266.05,    266.05,  266.05,  266.05,
  266,       266,     266,     266,
  265.85,    265.85,  265.85,  265.85,
  265.75,    265.75,  265.75,  265.75,
  265.85,    265.85,  265.85,  265.85,
  266.15,    266.15,  266.15,  266.15,
  266.55,    266.55,  266.55,  266.55,
  266.9,     266.9,   266.9,   266.9,
  267.15,    267.15,  267.15,  267.15,
  267.3,     267.3,   267.3,   267.3,
  267.45,    267.45,  267.45,  267.45,
  267.65,    267.65,  267.65,  267.65,
  267.85,    267.85,  267.85,  267.85,
  268.1,     268.1,   268.1,   268.1,
  268.35,    268.35,  268.35,  268.35,
  268.45,    268.45,  268.45,  268.45,
  268.5,     268.5,   268.5,   268.5,
  268.6,     268.6,   268.6,   268.6,
  268.75,    268.75,  268.75,  268.75,
  268.9,     268.9,   268.9,   268.9,
  269,       269,     269,     269,
  269.05,    269.05,  269.05,  269.05,
  269.1,     269.1,   269.1,   269.1,
  269.2,     269.2,   269.2,   269.2,
  269.25,    269.25,  269.25,  269.25,
  269.2,     269.2,   269.2,   269.2,
  269.15,    269.15,  269.15,  269.15,
  269.15,    269.15,  269.15,  269.15,
  269.15,    269.15,  269.15,  269.15,
  269.15,    269.15,  269.15,  269.15,
  269.1,     269.1,   269.1,   269.1,
  269,       269,     269,     269,
  268.95,    268.95,  268.95,  268.95,
  268.95,    268.95,  268.95,  268.95,
  268.9,     268.9,   268.9,   268.9,
  268.8,     268.8,   268.8,   268.8,
  268.8,     268.8,   268.8,   268.8,
  268.8,     268.8,   268.8,   268.8,
  268.75,    268.75,  268.75,  268.75,
  268.7,     268.7,   268.7,   268.7,
  268.65,    268.65,  268.65,  268.65,
  268.65,    268.65,  268.65,  268.65,
  268.75,    268.75,  268.75,  268.75,
  269,       269,     269,     269,
  269.2,     269.2,   269.2,   269.2,
  269.35,    269.35,  269.35,  269.35,
  269.5,     269.5,   269.5,   269.5,
  269.5,     269.5,   269.5,   269.5,
  269.45,    269.45,  269.45,  269.45,
  269.45,    269.45,  269.45,  269.45,
  269.45,    269.45,  269.45,  269.45,
  269.45,    269.45,  269.45,  269.45,
  269.4,     269.4,   269.4,   269.4,
  269.4,     269.4,   269.4,   269.4,
  269.45,    269.45,  269.45,  269.45,
  269.45,    269.45,  269.45,  269.45,
  269.5,     269.5,   269.5,   269.5,
  269.5,     269.5,   269.5,   269.5,
  269.5,     269.5,   269.5,   269.5,
  269.5,     269.5,   269.5,   269.5,
  269.5,     269.5,   269.5,   269.5,
  269.5,     269.5,   269.5,   269.5,
  269.5,     269.5,   269.5,   269.5,
  269.55,    269.55,  269.55,  269.55,
  269.55,    269.55,  269.55,  269.55,
  269.5,     269.5,   269.5,   269.5,
  269.45,    269.45,  269.45,  269.45,
  269.45,    269.45,  269.45,  269.45,
  269.4,     269.4,   269.4,   269.4,
  269.3,     269.3,   269.3,   269.3,
  269.3,     269.3,   269.3,   269.3,
  269.3,     269.3,   269.3,   269.3,
  269.2,     269.2,   269.2,   269.2,
  269.1,     269.1,   269.1,   269.1,
  269,       269,     269,     269,
  268.95,    268.95,  268.95,  268.95,
  268.95,    268.95,  268.95,  268.95,
  268.9,     268.9,   268.9,   268.9,
  268.85,    268.85,  268.85,  268.85,
  268.85,    268.85,  268.85,  268.85,
  268.8,     268.8,   268.8,   268.8,
  268.8,     268.8,   268.8,   268.8,
  268.85,    268.85,  268.85,  268.85,
  268.9,     268.9,   268.9,   268.9,
  269.05,    269.05,  269.05,  269.05,
  269.25,    269.25,  269.25,  269.25,
  269.45,    269.45,  269.45,  269.45,
  269.6,     269.6,   269.6,   269.6,
  269.65,    269.65,  269.65,  269.65,
  269.65,    269.65,  269.65,  269.65,
  269.65,    269.65,  269.65,  269.65,
  269.7,     269.7,   269.7,   269.7,
  269.8,     269.8,   269.8,   269.8,
  269.8,     269.8,   269.8,   269.8,
  269.8,     269.8,   269.8,   269.8,
  269.85,    269.85,  269.85,  269.85,
  269.85,    269.85,  269.85,  269.85,
  269.7,     269.7,   269.7,   269.7,
  269.5,     269.5,   269.5,   269.5,
  269.4,     269.4,   269.4,   269.4,
  269.3,     269.3,   269.3,   269.3,
  269.2,     269.2,   269.2,   269.2,
  269.1,     269.1,   269.1,   269.1,
  269,       269,     269,     269,
  268.8,     268.8,   268.8,   268.8,
  268.4,     268.4,   268.4,   268.4,
  267.95,    267.95,  267.95,  267.95,
  267.6,     267.6,   267.6,   267.6,
  267.3,     267.3,   267.3,   267.3,
  267,       267,     267,     267,
  266.85,    266.85,  266.85,  266.85,
  266.9,     266.9,   266.9,   266.9,
  267,       267,     267,     267,
  267.1,     267.1,   267.1,   267.1,
  267.05,    267.05,  267.05,  267.05,
  266.9,     266.9,   266.9,   266.9,
  266.85,    266.85,  266.85,  266.85,
  266.85,    266.85,  266.85,  266.85,
  266.8,     266.8,   266.8,   266.8,
  266.8,     266.8,   266.8,   266.8,
  267.05,    267.05,  267.05,  267.05,
  267.5,     267.5,   267.5,   267.5,
  267.9,     267.9,   267.9,   267.9,
  268.2,     268.2,   268.2,   268.2,
  268.5,     268.5,   268.5,   268.5,
  268.75,    268.75,  268.75,  268.75,
  268.9,     268.9,   268.9,   268.9,
  269,       269,     269,     269,
  269.1,     269.1,   269.1,   269.1,
  269.25,    269.25,  269.25,  269.25,
  269.4,     269.4,   269.4,   269.4,
  269.55,    269.55,  269.55,  269.55,
  269.75,    269.75,  269.75,  269.75,
  270.05,    270.05,  270.05,  270.05,
  270.55,    270.55,  270.55,  270.55,
  271.2,     271.2,   271.2,   271.2,
  271.8,     271.8,   271.8,   271.8,
  272.1,     272.1,   272.1,   272.1,
  272.35,    272.35,  272.35,  272.35,
  272.75,    272.75,  272.75,  272.75,
  273.15,    273.15,  273.15,  273.15,
  273.45,    273.45,  273.45,  273.45,
  273.6,     273.6,   273.6,   273.6,
  273.75,    273.75,  273.75,  273.75,
  273.95,    273.95,  273.95,  273.95,
  274.1,     274.1,   274.1,   274.1,
  274.15,    274.15,  274.15,  274.15,
  274.1,     274.1,   274.1,   274.1,
  274.1,     274.1,   274.1,   274.1,
  274.25,    274.25,  274.25,  274.25,
  274.4,     274.4,   274.4,   274.4,
  274.4,     274.4,   274.4,   274.4,
  274.4,     274.4,   274.4,   274.4,
  274.55,    274.55,  274.55,  274.55,
  274.65,    274.65,  274.65,  274.65,
  274.7,     274.7,   274.7,   274.7,
  274.7,     274.7,   274.7,   274.7,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.7,     274.7,   274.7,   274.7,
  274.75,    274.75,  274.75,  274.75,
  274.75,    274.75,  274.75,  274.75,
  274.75,    274.75,  274.75,  274.75,
  274.75,    274.75,  274.75,  274.75,
  274.8,     274.8,   274.8,   274.8,
  274.8,     274.8,   274.8,   274.8,
  274.7,     274.7,   274.7,   274.7,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.6,     274.6,   274.6,   274.6,
  274.5,     274.5,   274.5,   274.5,
  274.5,     274.5,   274.5,   274.5,
  274.55,    274.55,  274.55,  274.55,
  274.5,     274.5,   274.5,   274.5,
  274.45,    274.45,  274.45,  274.45,
  274.5,     274.5,   274.5,   274.5,
  274.6,     274.6,   274.6,   274.6,
  274.5,     274.5,   274.5,   274.5,
  274.5,     274.5,   274.5,   274.5,
  274.85,    274.85,  274.85,  274.85,
  275.55,    275.55,  275.55,  275.55,
  276.65,    276.65,  276.65,  276.65,
  277.65,    277.65,  277.65,  277.65,
  278.35,    278.35,  278.35,  278.35,
  278.95,    278.95,  278.95,  278.95,
  279.5,     279.5,   279.5,   279.5,
  279.9,     279.9,   279.9,   279.9,
  280.05,    280.05,  280.05,  280.05,
  280,       280,     280,     280,
  279.65,    279.65,  279.65,  279.65,
  278.95,    278.95,  278.95,  278.95,
  278.2,     278.2,   278.2,   278.2,
  277.6,     277.6,   277.6,   277.6,
  277.3,     277.3,   277.3,   277.3,
  276.9,     276.9,   276.9,   276.9,
  276.3,     276.3,   276.3,   276.3,
  275.85,    275.85,  275.85,  275.85,
  275.7,     275.7,   275.7,   275.7,
  275.7,     275.7,   275.7,   275.7,
  275.65,    275.65,  275.65,  275.65,
  275.4,     275.4,   275.4,   275.4,
  275,       275,     275,     275,
  274.75,    274.75,  274.75,  274.75,
  274.5,     274.5,   274.5,   274.5,
  274.25,    274.25,  274.25,  274.25,
  274.1,     274.1,   274.1,   274.1,
  274,       274,     274,     274,
  273.8,     273.8,   273.8,   273.8,
  273.6,     273.6,   273.6,   273.6,
  273.5,     273.5,   273.5,   273.5,
  273.4,     273.4,   273.4,   273.4,
  273.2,     273.2,   273.2,   273.2,
  273,       273,     273,     273,
  272.95,    272.95,  272.95,  272.95,
  272.9,     272.9,   272.9,   272.9,
  272.8,     272.8,   272.8,   272.8,
  272.65,    272.65,  272.65,  272.65,
  272.6,     272.6,   272.6,   272.6,
  272.75,    272.75,  272.75,  272.75,
  272.65,    272.65,  272.65,  272.65,
  272.35,    272.35,  272.35,  272.35,
  272.2,     272.2,   272.2,   272.2,
  272.15,    272.15,  272.15,  272.15,
  272.35,    272.35,  272.35,  272.35,
  273,       273,     273,     273,
  274.15,    274.15,  274.15,  274.15,
  275.85,    275.85,  275.85,  275.85,
  277.35,    277.35,  277.35,  277.35,
  278.3,     278.3,   278.3,   278.3,
  279.1,     279.1,   279.1,   279.1,
  280.1,     280.1,   280.1,   280.1,
  281.25,    281.25,  281.25,  281.25,
  282.1,     282.1,   282.1,   282.1,
  282.5,     282.5,   282.5,   282.5,
  282.55,    282.55,  282.55,  282.55,
  282.4,     282.4,   282.4,   282.4,
  282,       282,     282,     282,
  281.45,    281.45,  281.45,  281.45,
  280.6,     280.6,   280.6,   280.6,
  279.5,     279.5,   279.5,   279.5,
  278.5,     278.5,   278.5,   278.5,
  277.8,     277.8,   277.8,   277.8,
  277.45,    277.45,  277.45,  277.45,
  277.2,     277.2,   277.2,   277.2,
  276.75,    276.75,  276.75,  276.75,
  276.2,     276.2,   276.2,   276.2,
  275.55,    275.55,  275.55,  275.55,
  274.9,     274.9,   274.9,   274.9,
  274.55,    274.55,  274.55,  274.55,
  274.15,    274.15,  274.15,  274.15,
  273.65,    273.65,  273.65,  273.65,
  273.25,    273.25,  273.25,  273.25,
  273,       273,     273,     273,
  273.1,     273.1,   273.1,   273.1,
  273.3,     273.3,   273.3,   273.3,
  273.15,    273.15,  273.15,  273.15,
  272.8,     272.8,   272.8,   272.8,
  272.55,    272.55,  272.55,  272.55,
  272.3,     272.3,   272.3,   272.3,
  272,       272,     272,     272,
  271.7,     271.7,   271.7,   271.7,
  271.5,     271.5,   271.5,   271.5,
  271.35,    271.35,  271.35,  271.35,
  271.15,    271.15,  271.15,  271.15,
  270.95,    270.95,  270.95,  270.95,
  270.7,     270.7,   270.7,   270.7,
  270.5,     270.5,   270.5,   270.5,
  270.35,    270.35,  270.35,  270.35,
  270.2,     270.2,   270.2,   270.2,
  270.05,    270.05,  270.05,  270.05,
  269.9,     269.9,   269.9,   269.9,
  270,       270,     270,     270,
  270.35,    270.35,  270.35,  270.35,
  270.9,     270.9,   270.9,   270.9,
  271.8,     271.8,   271.8,   271.8,
  272.95,    272.95,  272.95,  272.95,
  274.05,    274.05,  274.05,  274.05,
  274.95,    274.95,  274.95,  274.95,
  275.65,    275.65,  275.65,  275.65,
  276.2,     276.2,   276.2,   276.2,
  276.75,    276.75,  276.75,  276.75,
  277.4,     277.4,   277.4,   277.4,
  277.8,     277.8,   277.8,   277.8,
  278.05,    278.05,  278.05,  278.05,
  278.2,     278.2,   278.2,   278.2,
  277.9,     277.9,   277.9,   277.9,
  277.2,     277.2,   277.2,   277.2,
  276.25,    276.25,  276.25,  276.25,
  275.65,    275.65,  275.65,  275.65,
  275.2,     275.2,   275.2,   275.2,
  274.5,     274.5,   274.5,   274.5,
  273.85,    273.85,  273.85,  273.85,
  273.45,    273.45,  273.45,  273.45,
  273.1,     273.1,   273.1,   273.1,
  272.7,     272.7,   272.7,   272.7,
  272.65,    272.65,  272.65,  272.65,
  272.6,     272.6,   272.6,   272.6,
  272.55,    272.55,  272.55,  272.55,
  272.55,    272.55,  272.55,  272.55,
  272.45,    272.45,  272.45,  272.45,
  272.35,    272.35,  272.35,  272.35,
  272.3,     272.3,   272.3,   272.3,
  272.3,     272.3,   272.3,   272.3,
  272.15,    272.15,  272.15,  272.15,
  271.65,    271.65,  271.65,  271.65,
  271.1,     271.1,   271.1,   271.1,
  270.95,    270.95,  270.95,  270.95,
  270.95,    270.95,  270.95,  270.95,
  270.85,    270.85,  270.85,  270.85,
  270.6,     270.6,   270.6,   270.6,
  270.35,    270.35,  270.35,  270.35,
  270.15,    270.15,  270.15,  270.15,
  269.9,     269.9,   269.9,   269.9,
  269.7,     269.7,   269.7,   269.7,
  269.7,     269.7,   269.7,   269.7,
  269.7,     269.7,   269.7,   269.7,
  269.6,     269.6,   269.6,   269.6,
  269.45,    269.45,  269.45,  269.45,
  269.35,    269.35,  269.35,  269.35,
  269.5,     269.5,   269.5,   269.5,
  270,       270,     270,     270,
  270.85,    270.85,  270.85,  270.85,
  272.05,    272.05,  272.05,  272.05,
  273.55,    273.55,  273.55,  273.55,
  275.1,     275.1,   275.1,   275.1,
  276.55,    276.55,  276.55,  276.55,
  277.8,     277.8,   277.8,   277.8,
  279,       279,     279,     279,
  279.85,    279.85,  279.85,  279.85,
  280.35,    280.35,  280.35,  280.35,
  280.9,     280.9,   280.9,   280.9,
  281.05,    281.05,  281.05,  281.05,
  280.95,    280.95,  280.95,  280.95,
  280.55,    280.55,  280.55,  280.55,
  279.3,     279.3,   279.3,   279.3,
  277.55,    277.55,  277.55,  277.55,
  276.25,    276.25,  276.25,  276.25,
  275.4,     275.4,   275.4,   275.4,
  274.65,    274.65,  274.65,  274.65,
  274.1,     274.1,   274.1,   274.1,
  273.7,     273.7,   273.7,   273.7,
  273.5,     273.5,   273.5,   273.5,
  273.4,     273.4,   273.4,   273.4,
  273.5,     273.5,   273.5,   273.5,
  273.6,     273.6,   273.6,   273.6,
  273.4,     273.4,   273.4,   273.4,
  273.2,     273.2,   273.2,   273.2,
  273.1,     273.1,   273.1,   273.1,
  273,       273,     273,     273,
  272.9,     272.9,   272.9,   272.9,
  272.75,    272.75,  272.75,  272.75,
  272.65,    272.65,  272.65,  272.65,
  272.4,     272.4,   272.4,   272.4,
  272.15,    272.15,  272.15,  272.15,
  272.2,     272.2,   272.2,   272.2,
  272.15,    272.15,  272.15,  272.15,
  272.2,     272.2,   272.2,   272.2,
  272.25,    272.25,  272.25,  272.25,
  272.3,     272.3,   272.3,   272.3,
  272.4,     272.4,   272.4,   272.4,
  272.25,    272.25,  272.25,  272.25,
  272.2,     272.2,   272.2,   272.2,
  272.35,    272.35,  272.35,  272.35,
  272.4,     272.4,   272.4,   272.4,
  272.2,     272.2,   272.2,   272.2,
  272,       272,     272,     272,
  272,       272,     272,     272,
  272.4,     272.4,   272.4,   272.4,
  273,       273,     273,     273,
  273.65,    273.65,  273.65,  273.65,
  274.7,     274.7,   274.7,   274.7,
  276.15,    276.15,  276.15,  276.15,
  277.55,    277.55,  277.55,  277.55,
  278.65,    278.65,  278.65,  278.65,
  279.45,    279.45,  279.45,  279.45,
  280,       280,     280,     280,
  280.5,     280.5,   280.5,   280.5,
  280.85,    280.85,  280.85,  280.85,
  281.05,    281.05,  281.05,  281.05,
  281.1,     281.1,   281.1,   281.1,
  280.95,    280.95,  280.95,  280.95,
  280.55,    280.55,  280.55,  280.55,
  279.9,     279.9,   279.9,   279.9,
  279.2,     279.2,   279.2,   279.2,
  278.55,    278.55,  278.55,  278.55,
  278.2,     278.2,   278.2,   278.2,
  278.15,    278.15,  278.15,  278.15,
  278.1,     278.1,   278.1,   278.1,
  278.05,    278.05,  278.05,  278.05,
  277.95,    277.95,  277.95,  277.95,
  277.8,     277.8,   277.8,   277.8,
  278,       278,     278,     278,
  278.5,     278.5,   278.5,   278.5,
  278.8,     278.8,   278.8,   278.8,
  278.95,    278.95,  278.95,  278.95,
  279,       279,     279,     279,
  278.85,    278.85,  278.85,  278.85,
  278.75,    278.75,  278.75,  278.75,
  278.75,    278.75,  278.75,  278.75,
  278.85,    278.85,  278.85,  278.85,
  278.8,     278.8,   278.8,   278.8,
  278.6,     278.6,   278.6,   278.6,
  278.5,     278.5,   278.5,   278.5,
  278.4,     278.4,   278.4,   278.4,
  278.2,     278.2,   278.2,   278.2,
  277.9,     277.9,   277.9,   277.9,
  277.65,    277.65,  277.65,  277.65,
  277.55,    277.55,  277.55,  277.55,
  277.55,    277.55,  277.55,  277.55,
  277.55,    277.55,  277.55,  277.55,
  277.55,    277.55,  277.55,  277.55,
  277.6,     277.6,   277.6,   277.6,
  277.65,    277.65,  277.65,  277.65,
  277.7,     277.7,   277.7,   277.7,
  277.85,    277.85,  277.85,  277.85,
  278,       278,     278,     278,
  278.1,     278.1,   278.1,   278.1,
  278.15,    278.15,  278.15,  278.15,
  278.2,     278.2,   278.2,   278.2,
  278.25,    278.25,  278.25,  278.25,
  278.2,     278.2,   278.2,   278.2,
  278.1,     278.1,   278.1,   278.1,
  278.05,    278.05,  278.05,  278.05,
  278.05,    278.05,  278.05,  278.05,
  278.05,    278.05,  278.05,  278.05,
  278.1,     278.1,   278.1,   278.1,
  278.1,     278.1,   278.1,   278.1,
  278.05,    278.05,  278.05,  278.05,
  277.95,    277.95,  277.95,  277.95,
  277.8,     277.8,   277.8,   277.8,
  277.7,     277.7,   277.7,   277.7,
  277.6,     277.6,   277.6,   277.6,
  277.5,     277.5,   277.5,   277.5,
  277.45,    277.45,  277.45,  277.45,
  277.4,     277.4,   277.4,   277.4,
  277.35,    277.35,  277.35,  277.35,
  277.3,     277.3,   277.3,   277.3,
  277.2,     277.2,   277.2,   277.2,
  277.1,     277.1,   277.1,   277.1,
  277,       277,     277,     277,
  276.9,     276.9,   276.9,   276.9,
  276.8,     276.8,   276.8,   276.8,
  276.75,    276.75,  276.75,  276.75,
  276.75,    276.75,  276.75,  276.75,
  276.75,    276.75,  276.75,  276.75,
  276.75,    276.75,  276.75,  276.75,
  276.65,    276.65,  276.65,  276.65,
  276.3,     276.3,   276.3,   276.3,
  275.6,     275.6,   275.6,   275.6,
  274.95,    274.95,  274.95,  274.95,
  274.65,    274.65,  274.65,  274.65,
  274.6,     274.6,   274.6,   274.6,
  274.8,     274.8,   274.8,   274.8,
  275.15,    275.15,  275.15,  275.15,
  275.45,    275.45,  275.45,  275.45,
  275.6,     275.6,   275.6,   275.6,
  275.7,     275.7,   275.7,   275.7,
  275.8,     275.8,   275.8,   275.8,
  275.9,     275.9,   275.9,   275.9,
  275.9,     275.9,   275.9,   275.9,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.9,     275.9,   275.9,   275.9,
  276,       276,     276,     276,
  276.15,    276.15,  276.15,  276.15,
  276.35,    276.35,  276.35,  276.35,
  276.5,     276.5,   276.5,   276.5,
  276.6,     276.6,   276.6,   276.6,
  276.6,     276.6,   276.6,   276.6,
  276.5,     276.5,   276.5,   276.5,
  276.45,    276.45,  276.45,  276.45,
  276.5,     276.5,   276.5,   276.5,
  276.55,    276.55,  276.55,  276.55,
  276.6,     276.6,   276.6,   276.6,
  276.75,    276.75,  276.75,  276.75,
  276.95,    276.95,  276.95,  276.95,
  277.05,    277.05,  277.05,  277.05,
  277.05,    277.05,  277.05,  277.05,
  277.05,    277.05,  277.05,  277.05,
  277,       277,     277,     277,
  276.95,    276.95,  276.95,  276.95,
  276.9,     276.9,   276.9,   276.9,
  276.9,     276.9,   276.9,   276.9,
  277,       277,     277,     277,
  277.1,     277.1,   277.1,   277.1,
  277.15,    277.15,  277.15,  277.15,
  277.15,    277.15,  277.15,  277.15,
  277.15,    277.15,  277.15,  277.15,
  277.1,     277.1,   277.1,   277.1,
  277,       277,     277,     277,
  276.9,     276.9,   276.9,   276.9,
  276.8,     276.8,   276.8,   276.8,
  276.7,     276.7,   276.7,   276.7,
  276.55,    276.55,  276.55,  276.55,
  276.4,     276.4,   276.4,   276.4,
  276.3,     276.3,   276.3,   276.3,
  276.2,     276.2,   276.2,   276.2,
  276.05,    276.05,  276.05,  276.05,
  275.65,    275.65,  275.65,  275.65,
  275.1,     275.1,   275.1,   275.1,
  274.75,    274.75,  274.75,  274.75,
  274.55,    274.55,  274.55,  274.55,
  274.4,     274.4,   274.4,   274.4,
  274.25,    274.25,  274.25,  274.25,
  274.05,    274.05,  274.05,  274.05,
  273.9,     273.9,   273.9,   273.9,
  273.9,     273.9,   273.9,   273.9,
  273.95,    273.95,  273.95,  273.95,
  274,       274,     274,     274,
  274.1,     274.1,   274.1,   274.1,
  274.15,    274.15,  274.15,  274.15,
  274.15,    274.15,  274.15,  274.15,
  274.2,     274.2,   274.2,   274.2,
  274.35,    274.35,  274.35,  274.35,
  274.55,    274.55,  274.55,  274.55,
  274.85,    274.85,  274.85,  274.85,
  275.25,    275.25,  275.25,  275.25,
  275.65,    275.65,  275.65,  275.65,
  276.1,     276.1,   276.1,   276.1,
  276.5,     276.5,   276.5,   276.5,
  276.7,     276.7,   276.7,   276.7,
  276.75,    276.75,  276.75,  276.75,
  276.8,     276.8,   276.8,   276.8,
  276.8,     276.8,   276.8,   276.8,
  276.65,    276.65,  276.65,  276.65,
  276.5,     276.5,   276.5,   276.5,
  276.35,    276.35,  276.35,  276.35,
  276.15,    276.15,  276.15,  276.15,
  276.05,    276.05,  276.05,  276.05,
  276.05,    276.05,  276.05,  276.05,
  276.05,    276.05,  276.05,  276.05,
  276,       276,     276,     276,
  275.9,     275.9,   275.9,   275.9,
  275.75,    275.75,  275.75,  275.75,
  275.5,     275.5,   275.5,   275.5,
  275.25,    275.25,  275.25,  275.25,
  275.05,    275.05,  275.05,  275.05,
  274.85,    274.85,  274.85,  274.85,
  274.45,    274.45,  274.45,  274.45,
  274.2,     274.2,   274.2,   274.2,
  274.25,    274.25,  274.25,  274.25,
  274.2,     274.2,   274.2,   274.2,
  274.1,     274.1,   274.1,   274.1,
  273.95,    273.95,  273.95,  273.95,
  273.9,     273.9,   273.9,   273.9,
  273.8,     273.8,   273.8,   273.8,
  273.55,    273.55,  273.55,  273.55,
  273.5,     273.5,   273.5,   273.5,
  273.65,    273.65,  273.65,  273.65,
  273.9,     273.9,   273.9,   273.9,
  274,       274,     274,     274,
  274,       274,     274,     274,
  274.05,    274.05,  274.05,  274.05,
  274.05,    274.05,  274.05,  274.05,
  274,       274,     274,     274,
  273.7,     273.7,   273.7,   273.7,
  273.3,     273.3,   273.3,   273.3,
  272.9,     272.9,   272.9,   272.9,
  272.6,     272.6,   272.6,   272.6,
  272.6,     272.6,   272.6,   272.6,
  272.8,     272.8,   272.8,   272.8,
  273,       273,     273,     273,
  273.3,     273.3,   273.3,   273.3,
  273.8,     273.8,   273.8,   273.8,
  274.15,    274.15,  274.15,  274.15,
  274.35,    274.35,  274.35,  274.35,
  274.6,     274.6,   274.6,   274.6,
  274.8,     274.8,   274.8,   274.8,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.8,     274.8,   274.8,   274.8,
  274.75,    274.75,  274.75,  274.75,
  274.7,     274.7,   274.7,   274.7,
  274.6,     274.6,   274.6,   274.6,
  274.55,    274.55,  274.55,  274.55,
  274.5,     274.5,   274.5,   274.5,
  274.3,     274.3,   274.3,   274.3,
  274,       274,     274,     274,
  273.85,    273.85,  273.85,  273.85,
  273.8,     273.8,   273.8,   273.8,
  273.85,    273.85,  273.85,  273.85,
  274,       274,     274,     274,
  273.95,    273.95,  273.95,  273.95,
  273.8,     273.8,   273.8,   273.8,
  273.6,     273.6,   273.6,   273.6,
  273.35,    273.35,  273.35,  273.35,
  273.1,     273.1,   273.1,   273.1,
  272.9,     272.9,   272.9,   272.9,
  272.8,     272.8,   272.8,   272.8,
  272.75,    272.75,  272.75,  272.75,
  272.75,    272.75,  272.75,  272.75,
  272.85,    272.85,  272.85,  272.85,
  273.05,    273.05,  273.05,  273.05,
  273.3,     273.3,   273.3,   273.3,
  273.5,     273.5,   273.5,   273.5,
  273.65,    273.65,  273.65,  273.65,
  273.8,     273.8,   273.8,   273.8,
  273.9,     273.9,   273.9,   273.9,
  273.95,    273.95,  273.95,  273.95,
  274.2,     274.2,   274.2,   274.2,
  274.7,     274.7,   274.7,   274.7,
  275.1,     275.1,   275.1,   275.1,
  275.35,    275.35,  275.35,  275.35,
  275.55,    275.55,  275.55,  275.55,
  275.75,    275.75,  275.75,  275.75,
  276,       276,     276,     276,
  276.25,    276.25,  276.25,  276.25,
  276.5,     276.5,   276.5,   276.5,
  276.8,     276.8,   276.8,   276.8,
  277.15,    277.15,  277.15,  277.15,
  277.8,     277.8,   277.8,   277.8,
  278.55,    278.55,  278.55,  278.55,
  279.15,    279.15,  279.15,  279.15,
  279.6,     279.6,   279.6,   279.6,
  280.05,    280.05,  280.05,  280.05,
  280.65,    280.65,  280.65,  280.65,
  281.45,    281.45,  281.45,  281.45,
  282.15,    282.15,  282.15,  282.15,
  282.2,     282.2,   282.2,   282.2,
  282.05,    282.05,  282.05,  282.05,
  281.9,     281.9,   281.9,   281.9,
  281.45,    281.45,  281.45,  281.45,
  280.95,    280.95,  280.95,  280.95,
  280.65,    280.65,  280.65,  280.65,
  280.55,    280.55,  280.55,  280.55,
  280.5,     280.5,   280.5,   280.5,
  280.5,     280.5,   280.5,   280.5,
  280.75,    280.75,  280.75,  280.75,
  280.85,    280.85,  280.85,  280.85,
  280.75,    280.75,  280.75,  280.75,
  280.55,    280.55,  280.55,  280.55,
  280.25,    280.25,  280.25,  280.25,
  280,       280,     280,     280,
  279.9,     279.9,   279.9,   279.9,
  280.1,     280.1,   280.1,   280.1,
  280.35,    280.35,  280.35,  280.35,
  280.35,    280.35,  280.35,  280.35,
  280.15,    280.15,  280.15,  280.15,
  279.65,    279.65,  279.65,  279.65,
  279,       279,     279,     279,
  278.85,    278.85,  278.85,  278.85,
  278.95,    278.95,  278.95,  278.95,
  278.65,    278.65,  278.65,  278.65,
  278.05,    278.05,  278.05,  278.05,
  277.6,     277.6,   277.6,   277.6,
  277.4,     277.4,   277.4,   277.4,
  277.4,     277.4,   277.4,   277.4,
  277.55,    277.55,  277.55,  277.55,
  277.65,    277.65,  277.65,  277.65,
  277.65,    277.65,  277.65,  277.65,
  277.75,    277.75,  277.75,  277.75,
  278,       278,     278,     278,
  278.2,     278.2,   278.2,   278.2,
  278.2,     278.2,   278.2,   278.2,
  278.2,     278.2,   278.2,   278.2,
  278.35,    278.35,  278.35,  278.35,
  278.6,     278.6,   278.6,   278.6,
  278.8,     278.8,   278.8,   278.8,
  278.95,    278.95,  278.95,  278.95,
  279.2,     279.2,   279.2,   279.2,
  279.6,     279.6,   279.6,   279.6,
  280,       280,     280,     280,
  280.2,     280.2,   280.2,   280.2,
  280.35,    280.35,  280.35,  280.35,
  280.45,    280.45,  280.45,  280.45,
  280.45,    280.45,  280.45,  280.45,
  280.55,    280.55,  280.55,  280.55,
  280.75,    280.75,  280.75,  280.75,
  280.55,    280.55,  280.55,  280.55,
  279.9,     279.9,   279.9,   279.9,
  279.15,    279.15,  279.15,  279.15,
  278.6,     278.6,   278.6,   278.6,
  278.3,     278.3,   278.3,   278.3,
  277.7,     277.7,   277.7,   277.7,
  277.05,    277.05,  277.05,  277.05,
  276.7,     276.7,   276.7,   276.7,
  276.5,     276.5,   276.5,   276.5,
  276.45,    276.45,  276.45,  276.45,
  276.3,     276.3,   276.3,   276.3,
  276.05,    276.05,  276.05,  276.05,
  275.9,     275.9,   275.9,   275.9,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  276.1,     276.1,   276.1,   276.1,
  276.5,     276.5,   276.5,   276.5,
  276.55,    276.55,  276.55,  276.55,
  276.7,     276.7,   276.7,   276.7,
  277.2,     277.2,   277.2,   277.2,
  277.2,     277.2,   277.2,   277.2,
  276.75,    276.75,  276.75,  276.75,
  276.8,     276.8,   276.8,   276.8,
  277.2,     277.2,   277.2,   277.2,
  277.1,     277.1,   277.1,   277.1,
  276.8,     276.8,   276.8,   276.8,
  276.8,     276.8,   276.8,   276.8,
  277,       277,     277,     277,
  277.2,     277.2,   277.2,   277.2,
  277.25,    277.25,  277.25,  277.25,
  277,       277,     277,     277,
  276.65,    276.65,  276.65,  276.65,
  276.5,     276.5,   276.5,   276.5,
  276.5,     276.5,   276.5,   276.5,
  276.55,    276.55,  276.55,  276.55,
  276.55,    276.55,  276.55,  276.55,
  276.3,     276.3,   276.3,   276.3,
  276.2,     276.2,   276.2,   276.2,
  276.75,    276.75,  276.75,  276.75,
  277.5,     277.5,   277.5,   277.5,
  277.85,    277.85,  277.85,  277.85,
  278.2,     278.2,   278.2,   278.2,
  278.85,    278.85,  278.85,  278.85,
  279.05,    279.05,  279.05,  279.05,
  278.85,    278.85,  278.85,  278.85,
  279.1,     279.1,   279.1,   279.1,
  279.4,     279.4,   279.4,   279.4,
  279.25,    279.25,  279.25,  279.25,
  278.9,     278.9,   278.9,   278.9,
  277.9,     277.9,   277.9,   277.9,
  276.8,     276.8,   276.8,   276.8,
  275.7,     275.7,   275.7,   275.7,
  274.6,     274.6,   274.6,   274.6,
  273.85,    273.85,  273.85,  273.85,
  273.4,     273.4,   273.4,   273.4,
  273.25,    273.25,  273.25,  273.25,
  272.85,    272.85,  272.85,  272.85,
  272.4,     272.4,   272.4,   272.4,
  272.3,     272.3,   272.3,   272.3,
  272.3,     272.3,   272.3,   272.3,
  272.2,     272.2,   272.2,   272.2,
  272,       272,     272,     272,
  271.75,    271.75,  271.75,  271.75,
  271.7,     271.7,   271.7,   271.7,
  271.5,     271.5,   271.5,   271.5,
  271.1,     271.1,   271.1,   271.1,
  271.1,     271.1,   271.1,   271.1,
  271.1,     271.1,   271.1,   271.1,
  271,       271,     271,     271,
  270.9,     270.9,   270.9,   270.9,
  270.85,    270.85,  270.85,  270.85,
  270.9,     270.9,   270.9,   270.9,
  270.7,     270.7,   270.7,   270.7,
  270.6,     270.6,   270.6,   270.6,
  270.65,    270.65,  270.65,  270.65,
  270.85,    270.85,  270.85,  270.85,
  270.75,    270.75,  270.75,  270.75,
  270.4,     270.4,   270.4,   270.4,
  270.45,    270.45,  270.45,  270.45,
  270.45,    270.45,  270.45,  270.45,
  270.45,    270.45,  270.45,  270.45,
  270.65,    270.65,  270.65,  270.65,
  271.05,    271.05,  271.05,  271.05,
  271.5,     271.5,   271.5,   271.5,
  272.1,     272.1,   272.1,   272.1,
  273.1,     273.1,   273.1,   273.1,
  274.45,    274.45,  274.45,  274.45,
  276,       276,     276,     276,
  277.5,     277.5,   277.5,   277.5,
  278.5,     278.5,   278.5,   278.5,
  279.25,    279.25,  279.25,  279.25,
  280,       280,     280,     280,
  280.2,     280.2,   280.2,   280.2,
  280.25,    280.25,  280.25,  280.25,
  280,       280,     280,     280,
  279.45,    279.45,  279.45,  279.45,
  278.95,    278.95,  278.95,  278.95,
  278.05,    278.05,  278.05,  278.05,
  275.95,    275.95,  275.95,  275.95,
  273.6,     273.6,   273.6,   273.6,
  272.4,     272.4,   272.4,   272.4,
  272,       272,     272,     272,
  272,       272,     272,     272,
  271.95,    271.95,  271.95,  271.95,
  271.95,    271.95,  271.95,  271.95,
  272.15,    272.15,  272.15,  272.15,
  272.3,     272.3,   272.3,   272.3,
  272.35,    272.35,  272.35,  272.35,
  272.35,    272.35,  272.35,  272.35,
  272.4,     272.4,   272.4,   272.4,
  272.5,     272.5,   272.5,   272.5,
  272.55,    272.55,  272.55,  272.55,
  272.5,     272.5,   272.5,   272.5,
  272.5,     272.5,   272.5,   272.5,
  272.7,     272.7,   272.7,   272.7,
  272.9,     272.9,   272.9,   272.9,
  272.95,    272.95,  272.95,  272.95,
  272.95,    272.95,  272.95,  272.95,
  273,       273,     273,     273,
  273,       273,     273,     273,
  272.95,    272.95,  272.95,  272.95,
  273,       273,     273,     273,
  273.1,     273.1,   273.1,   273.1,
  273.2,     273.2,   273.2,   273.2,
  273.3,     273.3,   273.3,   273.3,
  273.45,    273.45,  273.45,  273.45,
  273.55,    273.55,  273.55,  273.55,
  273.65,    273.65,  273.65,  273.65,
  273.8,     273.8,   273.8,   273.8,
  273.75,    273.75,  273.75,  273.75,
  273.55,    273.55,  273.55,  273.55,
  273.4,     273.4,   273.4,   273.4,
  273.35,    273.35,  273.35,  273.35,
  273.3,     273.3,   273.3,   273.3,
  273.25,    273.25,  273.25,  273.25,
  273.25,    273.25,  273.25,  273.25,
  273.2,     273.2,   273.2,   273.2,
  273.15,    273.15,  273.15,  273.15,
  273.15,    273.15,  273.15,  273.15,
  273.2,     273.2,   273.2,   273.2,
  273.15,    273.15,  273.15,  273.15,
  273,       273,     273,     273,
  272.85,    272.85,  272.85,  272.85,
  272.65,    272.65,  272.65,  272.65,
  272.45,    272.45,  272.45,  272.45,
  272.3,     272.3,   272.3,   272.3,
  272.25,    272.25,  272.25,  272.25,
  272.2,     272.2,   272.2,   272.2,
  272.2,     272.2,   272.2,   272.2,
  272.1,     272.1,   272.1,   272.1,
  271.8,     271.8,   271.8,   271.8,
  271.5,     271.5,   271.5,   271.5,
  271.25,    271.25,  271.25,  271.25,
  271,       271,     271,     271,
  270.75,    270.75,  270.75,  270.75,
  270.65,    270.65,  270.65,  270.65,
  270.5,     270.5,   270.5,   270.5,
  270.25,    270.25,  270.25,  270.25,
  270,       270,     270,     270,
  269.75,    269.75,  269.75,  269.75,
  269.55,    269.55,  269.55,  269.55,
  269.35,    269.35,  269.35,  269.35,
  269.2,     269.2,   269.2,   269.2,
  269.1,     269.1,   269.1,   269.1,
  269,       269,     269,     269,
  268.85,    268.85,  268.85,  268.85,
  268.65,    268.65,  268.65,  268.65,
  268.65,    268.65,  268.65,  268.65,
  268.85,    268.85,  268.85,  268.85,
  268.95,    268.95,  268.95,  268.95,
  268.9,     268.9,   268.9,   268.9,
  268.85,    268.85,  268.85,  268.85,
  268.8,     268.8,   268.8,   268.8,
  268.65,    268.65,  268.65,  268.65,
  268.4,     268.4,   268.4,   268.4,
  268.2,     268.2,   268.2,   268.2,
  268.05,    268.05,  268.05,  268.05,
  267.75,    267.75,  267.75,  267.75,
  267.7,     267.7,   267.7,   267.7,
  268,       268,     268,     268,
  268.2,     268.2,   268.2,   268.2,
  268.55,    268.55,  268.55,  268.55,
  269.15,    269.15,  269.15,  269.15,
  269.75,    269.75,  269.75,  269.75,
  270.25,    270.25,  270.25,  270.25,
  270.65,    270.65,  270.65,  270.65,
  271.1,     271.1,   271.1,   271.1,
  271.35,    271.35,  271.35,  271.35,
  271.45,    271.45,  271.45,  271.45,
  271.65,    271.65,  271.65,  271.65,
  271.75,    271.75,  271.75,  271.75,
  271.75,    271.75,  271.75,  271.75,
  271.75,    271.75,  271.75,  271.75,
  271.75,    271.75,  271.75,  271.75,
  271.65,    271.65,  271.65,  271.65,
  271.4,     271.4,   271.4,   271.4,
  271.25,    271.25,  271.25,  271.25,
  271.2,     271.2,   271.2,   271.2,
  271.1,     271.1,   271.1,   271.1,
  270.9,     270.9,   270.9,   270.9,
  270.8,     270.8,   270.8,   270.8,
  270.7,     270.7,   270.7,   270.7,
  270.35,    270.35,  270.35,  270.35,
  269.85,    269.85,  269.85,  269.85,
  269.65,    269.65,  269.65,  269.65,
  270,       270,     270,     270,
  270.05,    270.05,  270.05,  270.05,
  269.55,    269.55,  269.55,  269.55,
  269.15,    269.15,  269.15,  269.15,
  269.2,     269.2,   269.2,   269.2,
  269.45,    269.45,  269.45,  269.45,
  269.7,     269.7,   269.7,   269.7,
  270,       270,     270,     270,
  270.3,     270.3,   270.3,   270.3,
  270.6,     270.6,   270.6,   270.6,
  270.95,    270.95,  270.95,  270.95,
  271.25,    271.25,  271.25,  271.25,
  271.45,    271.45,  271.45,  271.45,
  271.55,    271.55,  271.55,  271.55,
  271.8,     271.8,   271.8,   271.8,
  272.15,    272.15,  272.15,  272.15,
  272.4,     272.4,   272.4,   272.4,
  272.65,    272.65,  272.65,  272.65,
  272.9,     272.9,   272.9,   272.9,
  273.15,    273.15,  273.15,  273.15,
  273.3,     273.3,   273.3,   273.3,
  273.35,    273.35,  273.35,  273.35,
  273.45,    273.45,  273.45,  273.45,
  273.65,    273.65,  273.65,  273.65,
  274,       274,     274,     274,
  274.45,    274.45,  274.45,  274.45,
  274.9,     274.9,   274.9,   274.9,
  275.25,    275.25,  275.25,  275.25,
  275.5,     275.5,   275.5,   275.5,
  275.75,    275.75,  275.75,  275.75,
  275.95,    275.95,  275.95,  275.95,
  276.05,    276.05,  276.05,  276.05,
  275.95,    275.95,  275.95,  275.95,
  275.8,     275.8,   275.8,   275.8,
  275.75,    275.75,  275.75,  275.75,
  275.75,    275.75,  275.75,  275.75,
  275.8,     275.8,   275.8,   275.8,
  275.75,    275.75,  275.75,  275.75,
  275.6,     275.6,   275.6,   275.6,
  275.6,     275.6,   275.6,   275.6,
  275.65,    275.65,  275.65,  275.65,
  275.65,    275.65,  275.65,  275.65,
  275.65,    275.65,  275.65,  275.65,
  275.7,     275.7,   275.7,   275.7,
  275.7,     275.7,   275.7,   275.7,
  275.7,     275.7,   275.7,   275.7,
  275.8,     275.8,   275.8,   275.8,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.75,    275.75,  275.75,  275.75,
  275.6,     275.6,   275.6,   275.6,
  275.5,     275.5,   275.5,   275.5,
  275.4,     275.4,   275.4,   275.4,
  275.3,     275.3,   275.3,   275.3,
  275.2,     275.2,   275.2,   275.2,
  275.15,    275.15,  275.15,  275.15,
  275.2,     275.2,   275.2,   275.2,
  275.3,     275.3,   275.3,   275.3,
  275.35,    275.35,  275.35,  275.35,
  275.35,    275.35,  275.35,  275.35,
  275.35,    275.35,  275.35,  275.35,
  275.3,     275.3,   275.3,   275.3,
  275.25,    275.25,  275.25,  275.25,
  275.2,     275.2,   275.2,   275.2,
  275.05,    275.05,  275.05,  275.05,
  274.8,     274.8,   274.8,   274.8,
  274.55,    274.55,  274.55,  274.55,
  274.45,    274.45,  274.45,  274.45,
  274.5,     274.5,   274.5,   274.5,
  274.65,    274.65,  274.65,  274.65,
  274.8,     274.8,   274.8,   274.8,
  274.95,    274.95,  274.95,  274.95,
  275.05,    275.05,  275.05,  275.05,
  275.1,     275.1,   275.1,   275.1,
  275.2,     275.2,   275.2,   275.2,
  275.35,    275.35,  275.35,  275.35,
  275.5,     275.5,   275.5,   275.5,
  275.5,     275.5,   275.5,   275.5,
  275.45,    275.45,  275.45,  275.45,
  275.45,    275.45,  275.45,  275.45,
  275.45,    275.45,  275.45,  275.45,
  275.45,    275.45,  275.45,  275.45,
  275.4,     275.4,   275.4,   275.4,
  275.35,    275.35,  275.35,  275.35,
  275.35,    275.35,  275.35,  275.35,
  275.3,     275.3,   275.3,   275.3,
  275.25,    275.25,  275.25,  275.25,
  275.2,     275.2,   275.2,   275.2,
  275.1,     275.1,   275.1,   275.1,
  275,       275,     275,     275,
  274.9,     274.9,   274.9,   274.9,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.8,     274.8,   274.8,   274.8,
  274.75,    274.75,  274.75,  274.75,
  274.75,    274.75,  274.75,  274.75,
  274.75,    274.75,  274.75,  274.75,
  274.7,     274.7,   274.7,   274.7,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.6,     274.6,   274.6,   274.6,
  274.4,     274.4,   274.4,   274.4,
  274.25,    274.25,  274.25,  274.25,
  274.35,    274.35,  274.35,  274.35,
  274.3,     274.3,   274.3,   274.3,
  274.1,     274.1,   274.1,   274.1,
  274.05,    274.05,  274.05,  274.05,
  274.2,     274.2,   274.2,   274.2,
  274.4,     274.4,   274.4,   274.4,
  274.55,    274.55,  274.55,  274.55,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.85,    274.85,  274.85,  274.85,
  275.05,    275.05,  275.05,  275.05,
  275.05,    275.05,  275.05,  275.05,
  275.1,     275.1,   275.1,   275.1,
  275.25,    275.25,  275.25,  275.25,
  275.45,    275.45,  275.45,  275.45,
  275.55,    275.55,  275.55,  275.55,
  275.6,     275.6,   275.6,   275.6,
  275.7,     275.7,   275.7,   275.7,
  275.8,     275.8,   275.8,   275.8,
  275.9,     275.9,   275.9,   275.9,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.95,    275.95,  275.95,  275.95,
  275.9,     275.9,   275.9,   275.9,
  275.8,     275.8,   275.8,   275.8,
  275.7,     275.7,   275.7,   275.7,
  275.65,    275.65,  275.65,  275.65,
  275.65,    275.65,  275.65,  275.65,
  275.65,    275.65,  275.65,  275.65,
  275.6,     275.6,   275.6,   275.6,
  275.5,     275.5,   275.5,   275.5,
  275.4,     275.4,   275.4,   275.4,
  275.35,    275.35,  275.35,  275.35,
  275.35,    275.35,  275.35,  275.35,
  275.3,     275.3,   275.3,   275.3,
  275.25,    275.25,  275.25,  275.25,
  275.2,     275.2,   275.2,   275.2,
  275.15,    275.15,  275.15,  275.15,
  275.15,    275.15,  275.15,  275.15,
  275.15,    275.15,  275.15,  275.15,
  275.1,     275.1,   275.1,   275.1,
  275.05,    275.05,  275.05,  275.05,
  275,       275,     275,     275,
  275,       275,     275,     275,
  275,       275,     275,     275,
  274.95,    274.95,  274.95,  274.95,
  274.95,    274.95,  274.95,  274.95,
  274.9,     274.9,   274.9,   274.9,
  274.65,    274.65,  274.65,  274.65,
  274.2,     274.2,   274.2,   274.2,
  273.85,    273.85,  273.85,  273.85,
  273.6,     273.6,   273.6,   273.6,
  273.35,    273.35,  273.35,  273.35,
  273.1,     273.1,   273.1,   273.1,
  273,       273,     273,     273,
  273.3,     273.3,   273.3,   273.3,
  273.65,    273.65,  273.65,  273.65,
  273.85,    273.85,  273.85,  273.85,
  274.1,     274.1,   274.1,   274.1,
  274.4,     274.4,   274.4,   274.4,
  274.7,     274.7,   274.7,   274.7,
  275,       275,     275,     275,
  275.25,    275.25,  275.25,  275.25,
  275.5,     275.5,   275.5,   275.5,
  275.9,     275.9,   275.9,   275.9,
  276.3,     276.3,   276.3,   276.3,
  276.5,     276.5,   276.5,   276.5,
  276.5,     276.5,   276.5,   276.5,
  276.35,    276.35,  276.35,  276.35,
  276.3,     276.3,   276.3,   276.3,
  276.55,    276.55,  276.55,  276.55,
  276.75,    276.75,  276.75,  276.75,
  276.7,     276.7,   276.7,   276.7,
  276.45,    276.45,  276.45,  276.45,
  276.15,    276.15,  276.15,  276.15,
  275.95,    275.95,  275.95,  275.95,
  275.75,    275.75,  275.75,  275.75,
  275.5,     275.5,   275.5,   275.5,
  275.3,     275.3,   275.3,   275.3,
  275.25,    275.25,  275.25,  275.25,
  275.25,    275.25,  275.25,  275.25,
  275.2,     275.2,   275.2,   275.2,
  275.15,    275.15,  275.15,  275.15,
  275.1,     275.1,   275.1,   275.1,
  275.1,     275.1,   275.1,   275.1,
  275.1,     275.1,   275.1,   275.1,
  275,       275,     275,     275,
  274.9,     274.9,   274.9,   274.9,
  274.85,    274.85,  274.85,  274.85,
  274.75,    274.75,  274.75,  274.75,
  274.65,    274.65,  274.65,  274.65,
  274.45,    274.45,  274.45,  274.45,
  274.35,    274.35,  274.35,  274.35,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.5,     274.5,   274.5,   274.5,
  274.55,    274.55,  274.55,  274.55,
  274.6,     274.6,   274.6,   274.6,
  274.7,     274.7,   274.7,   274.7,
  274.7,     274.7,   274.7,   274.7,
  274.55,    274.55,  274.55,  274.55,
  274.5,     274.5,   274.5,   274.5,
  274.45,    274.45,  274.45,  274.45,
  274.35,    274.35,  274.35,  274.35,
  274.3,     274.3,   274.3,   274.3,
  274.3,     274.3,   274.3,   274.3,
  274.3,     274.3,   274.3,   274.3,
  274.3,     274.3,   274.3,   274.3,
  274.5,     274.5,   274.5,   274.5,
  274.7,     274.7,   274.7,   274.7,
  274.85,    274.85,  274.85,  274.85,
  275,       275,     275,     275,
  275.15,    275.15,  275.15,  275.15,
  275.25,    275.25,  275.25,  275.25,
  275.3,     275.3,   275.3,   275.3,
  275.35,    275.35,  275.35,  275.35,
  275.4,     275.4,   275.4,   275.4,
  275.35,    275.35,  275.35,  275.35,
  275.25,    275.25,  275.25,  275.25,
  275.15,    275.15,  275.15,  275.15,
  275,       275,     275,     275,
  274.85,    274.85,  274.85,  274.85,
  274.7,     274.7,   274.7,   274.7,
  274.55,    274.55,  274.55,  274.55,
  274.3,     274.3,   274.3,   274.3,
  273.9,     273.9,   273.9,   273.9,
  273.6,     273.6,   273.6,   273.6,
  273.6,     273.6,   273.6,   273.6,
  273.65,    273.65,  273.65,  273.65,
  273.35,    273.35,  273.35,  273.35,
  272.75,    272.75,  272.75,  272.75,
  272.25,    272.25,  272.25,  272.25,
  271.9,     271.9,   271.9,   271.9,
  271.8,     271.8,   271.8,   271.8,
  271.85,    271.85,  271.85,  271.85,
  271.8,     271.8,   271.8,   271.8,
  271.7,     271.7,   271.7,   271.7,
  271.55,    271.55,  271.55,  271.55,
  271.45,    271.45,  271.45,  271.45,
  271.35,    271.35,  271.35,  271.35,
  271.25,    271.25,  271.25,  271.25,
  271.25,    271.25,  271.25,  271.25,
  271.1,     271.1,   271.1,   271.1,
  270.85,    270.85,  270.85,  270.85,
  270.7,     270.7,   270.7,   270.7,
  270.6,     270.6,   270.6,   270.6,
  270.5,     270.5,   270.5,   270.5,
  270.4,     270.4,   270.4,   270.4,
  270.3,     270.3,   270.3,   270.3,
  270.35,    270.35,  270.35,  270.35,
  270.4,     270.4,   270.4,   270.4,
  270.4,     270.4,   270.4,   270.4,
  270.45,    270.45,  270.45,  270.45,
  270.5,     270.5,   270.5,   270.5,
  270.85,    270.85,  270.85,  270.85,
  271.6,     271.6,   271.6,   271.6,
  272.45,    272.45,  272.45,  272.45,
  273.35,    273.35,  273.35,  273.35,
  273.9,     273.9,   273.9,   273.9,
  274,       274,     274,     274,
  274.15,    274.15,  274.15,  274.15,
  274.55,    274.55,  274.55,  274.55,
  274.85,    274.85,  274.85,  274.85,
  274.4,     274.4,   274.4,   274.4,
  273.9,     273.9,   273.9,   273.9,
  273.7,     273.7,   273.7,   273.7,
  273.35,    273.35,  273.35,  273.35,
  273.1,     273.1,   273.1,   273.1,
  273.05,    273.05,  273.05,  273.05,
  273,       273,     273,     273,
  273,       273,     273,     273,
  273,       273,     273,     273,
  272.95,    272.95,  272.95,  272.95,
  273,       273,     273,     273,
  273.05,    273.05,  273.05,  273.05,
  273.1,     273.1,   273.1,   273.1,
  273.2,     273.2,   273.2,   273.2,
  273.3,     273.3,   273.3,   273.3,
  273.35,    273.35,  273.35,  273.35,
  273.4,     273.4,   273.4,   273.4,
  273.45,    273.45,  273.45,  273.45,
  273.5,     273.5,   273.5,   273.5,
  273.55,    273.55,  273.55,  273.55,
  273.55,    273.55,  273.55,  273.55,
  273.6,     273.6,   273.6,   273.6,
  273.65,    273.65,  273.65,  273.65,
  273.7,     273.7,   273.7,   273.7,
  273.75,    273.75,  273.75,  273.75,
  273.75,    273.75,  273.75,  273.75,
  273.75,    273.75,  273.75,  273.75,
  273.75,    273.75,  273.75,  273.75,
  273.75,    273.75,  273.75,  273.75,
  273.75,    273.75,  273.75,  273.75,
  273.85,    273.85,  273.85,  273.85,
  274,       274,     274,     274,
  274,       274,     274,     274,
  273.9,     273.9,   273.9,   273.9,
  273.7,     273.7,   273.7,   273.7,
  273.55,    273.55,  273.55,  273.55,
  273.5,     273.5,   273.5,   273.5,
  273.4,     273.4,   273.4,   273.4,
  273.35,    273.35,  273.35,  273.35,
  273.4,     273.4,   273.4,   273.4,
  273.55,    273.55,  273.55,  273.55,
  273.8,     273.8,   273.8,   273.8,
  274,       274,     274,     274,
  274.1,     274.1,   274.1,   274.1,
  274.15,    274.15,  274.15,  274.15,
  274.25,    274.25,  274.25,  274.25,
  274.4,     274.4,   274.4,   274.4,
  274.3,     274.3,   274.3,   274.3,
  273.95,    273.95,  273.95,  273.95,
  273.75,    273.75,  273.75,  273.75,
  273.75,    273.75,  273.75,  273.75,
  273.8,     273.8,   273.8,   273.8,
  273.9,     273.9,   273.9,   273.9,
  274.1,     274.1,   274.1,   274.1,
  274.3,     274.3,   274.3,   274.3,
  274.35,    274.35,  274.35,  274.35,
  274.3,     274.3,   274.3,   274.3,
  274.1,     274.1,   274.1,   274.1,
  273.95,    273.95,  273.95,  273.95,
  273.95,    273.95,  273.95,  273.95,
  273.95,    273.95,  273.95,  273.95,
  273.8,     273.8,   273.8,   273.8,
  273.6,     273.6,   273.6,   273.6,
  273.5,     273.5,   273.5,   273.5,
  273.55,    273.55,  273.55,  273.55,
  273.75,    273.75,  273.75,  273.75,
  273.95,    273.95,  273.95,  273.95,
  274.15,    274.15,  274.15,  274.15,
  274.2,     274.2,   274.2,   274.2,
  274.05,    274.05,  274.05,  274.05,
  273.8,     273.8,   273.8,   273.8,
  273.55,    273.55,  273.55,  273.55,
  273.45,    273.45,  273.45,  273.45,
  273.45,    273.45,  273.45,  273.45,
  273.45,    273.45,  273.45,  273.45,
  273.5,     273.5,   273.5,   273.5,
  273.65,    273.65,  273.65,  273.65,
  273.85,    273.85,  273.85,  273.85,
  274.1,     274.1,   274.1,   274.1,
  274.4,     274.4,   274.4,   274.4,
  274.7,     274.7,   274.7,   274.7,
  274.95,    274.95,  274.95,  274.95,
  275.15,    275.15,  275.15,  275.15,
  275.25,    275.25,  275.25,  275.25,
  275.3,     275.3,   275.3,   275.3,
  275.4,     275.4,   275.4,   275.4,
  275.6,     275.6,   275.6,   275.6,
  275.95,    275.95,  275.95,  275.95,
  276.25,    276.25,  276.25,  276.25,
  276.45,    276.45,  276.45,  276.45,
  276.75,    276.75,  276.75,  276.75,
  277.1,     277.1,   277.1,   277.1,
  277.3,     277.3,   277.3,   277.3,
  277.4,     277.4,   277.4,   277.4,
  277.5,     277.5,   277.5,   277.5,
  277.65,    277.65,  277.65,  277.65,
  277.85,    277.85,  277.85,  277.85,
  278.05,    278.05,  278.05,  278.05,
  278.15,    278.15,  278.15,  278.15,
  278.15,    278.15,  278.15,  278.15,
  278.25,    278.25,  278.25,  278.25,
  278.4,     278.4,   278.4,   278.4,
  278.55,    278.55,  278.55,  278.55,
  278.75,    278.75,  278.75,  278.75,
  278.9,     278.9,   278.9,   278.9,
  279,       279,     279,     279,
  279.05,    279.05,  279.05,  279.05,
  279.05,    279.05,  279.05,  279.05,
  279.05,    279.05,  279.05,  279.05,
  279.15,    279.15,  279.15,  279.15,
  279.25,    279.25,  279.25,  279.25,
  279.3,     279.3,   279.3,   279.3,
  279.4,     279.4,   279.4,   279.4,
  279.4,     279.4,   279.4,   279.4,
  279.35,    279.35,  279.35,  279.35,
  279.3,     279.3,   279.3,   279.3,
  279.2,     279.2,   279.2,   279.2,
  279.15,    279.15,  279.15,  279.15,
  279.05,    279.05,  279.05,  279.05,
  278.2,     278.2,   278.2,   278.2,
  276.9,     276.9,   276.9,   276.9,
  276.25,    276.25,  276.25,  276.25,
  276.15,    276.15,  276.15,  276.15,
  276.1,     276.1,   276.1,   276.1,
  276,       276,     276,     276,
  275.9,     275.9,   275.9,   275.9,
  275.9,     275.9,   275.9,   275.9,
  275.9,     275.9,   275.9,   275.9,
  275.85,    275.85,  275.85,  275.85,
  275.8,     275.8,   275.8,   275.8,
  275.65,    275.65,  275.65,  275.65,
  275.45,    275.45,  275.45,  275.45,
  275.25,    275.25,  275.25,  275.25,
  275.2,     275.2,   275.2,   275.2,
  275.2,     275.2,   275.2,   275.2,
  275,       275,     275,     275,
  275.1,     275.1,   275.1,   275.1,
  275.8,     275.8,   275.8,   275.8,
  276.6,     276.6,   276.6,   276.6,
  277.2,     277.2,   277.2,   277.2,
  277.7,     277.7,   277.7,   277.7,
  278.15,    278.15,  278.15,  278.15,
  278.4,     278.4,   278.4,   278.4,
  278.6,     278.6,   278.6,   278.6,
  278.65,    278.65,  278.65,  278.65,
  278.45,    278.45,  278.45,  278.45,
  278.35,    278.35,  278.35,  278.35,
  278.4,     278.4,   278.4,   278.4,
  278.3,     278.3,   278.3,   278.3,
  278.1,     278.1,   278.1,   278.1,
  277.95,    277.95,  277.95,  277.95,
  277.65,    277.65,  277.65,  277.65,
  277.1,     277.1,   277.1,   277.1,
  276.45,    276.45,  276.45,  276.45,
  275.9,     275.9,   275.9,   275.9,
  275.5,     275.5,   275.5,   275.5,
  275.35,    275.35,  275.35,  275.35,
  275.4,     275.4,   275.4,   275.4,
  275.25,    275.25,  275.25,  275.25,
  274.8,     274.8,   274.8,   274.8,
  274.4,     274.4,   274.4,   274.4,
  274.2,     274.2,   274.2,   274.2,
  274.15,    274.15,  274.15,  274.15,
  274.1,     274.1,   274.1,   274.1,
  274.05,    274.05,  274.05,  274.05,
  274.1,     274.1,   274.1,   274.1,
  274.2,     274.2,   274.2,   274.2,
  274.25,    274.25,  274.25,  274.25,
  274.35,    274.35,  274.35,  274.35,
  274.45,    274.45,  274.45,  274.45,
  274.5,     274.5,   274.5,   274.5,
  274.65,    274.65,  274.65,  274.65,
  274.85,    274.85,  274.85,  274.85,
  275,       275,     275,     275,
  275.05,    275.05,  275.05,  275.05,
  275,       275,     275,     275,
  274.95,    274.95,  274.95,  274.95,
  274.85,    274.85,  274.85,  274.85,
  274.7,     274.7,   274.7,   274.7,
  274.6,     274.6,   274.6,   274.6,
  274.55,    274.55,  274.55,  274.55,
  274.55,    274.55,  274.55,  274.55,
  274.55,    274.55,  274.55,  274.55,
  274.65,    274.65,  274.65,  274.65,
  274.9,     274.9,   274.9,   274.9,
  275.2,     275.2,   275.2,   275.2,
  275.55,    275.55,  275.55,  275.55,
  276,       276,     276,     276,
  276.65,    276.65,  276.65,  276.65,
  277.5,     277.5,   277.5,   277.5,
  278.35,    278.35,  278.35,  278.35,
  279.1,     279.1,   279.1,   279.1,
  279.7,     279.7,   279.7,   279.7,
  280.1,     280.1,   280.1,   280.1,
  280.3,     280.3,   280.3,   280.3,
  280.35,    280.35,  280.35,  280.35,
  280.45,    280.45,  280.45,  280.45,
  280.6,     280.6,   280.6,   280.6,
  280.65,    280.65,  280.65,  280.65,
  280.65,    280.65,  280.65,  280.65,
  280.65,    280.65,  280.65,  280.65,
  280.55,    280.55,  280.55,  280.55,
  280.35,    280.35,  280.35,  280.35,
  280.1,     280.1,   280.1,   280.1,
  279.75,    279.75,  279.75,  279.75,
  279.25,    279.25,  279.25,  279.25,
  278.8,     278.8,   278.8,   278.8,
  278.5,     278.5,   278.5,   278.5,
  278.25,    278.25,  278.25,  278.25,
  278.15,    278.15,  278.15,  278.15,
  278.05,    278.05,  278.05,  278.05,
  277.85,    277.85,  277.85,  277.85,
  277.85,    277.85,  277.85,  277.85,
  277.95,    277.95,  277.95,  277.95,
  277.9,     277.9,   277.9,   277.9,
  277.8,     277.8,   277.8,   277.8,
  277.65,    277.65,  277.65,  277.65,
  277.55,    277.55,  277.55,  277.55,
  277.5,     277.5,   277.5,   277.5,
  277.55,    277.55,  277.55,  277.55,
  277.75,    277.75,  277.75,  277.75,
  277.9,     277.9,   277.9,   277.9,
  277.95,    277.95,  277.95,  277.95,
  278,       278,     278,     278,
  278.1,     278.1,   278.1,   278.1,
  278.15,    278.15,  278.15,  278.15,
  278.15,    278.15,  278.15,  278.15,
  278.2,     278.2,   278.2,   278.2,
  278.3,     278.3,   278.3,   278.3,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.4,     278.4,   278.4,   278.4,
  278.65,    278.65,  278.65,  278.65,
  279.2,     279.2,   279.2,   279.2,
  279.75,    279.75,  279.75,  279.75,
  280.15,    280.15,  280.15,  280.15,
  280.4,     280.4,   280.4,   280.4,
  280.7,     280.7,   280.7,   280.7,
  281.55,    281.55,  281.55,  281.55,
  282.25,    282.25,  282.25,  282.25,
  282.25,    282.25,  282.25,  282.25,
  282.05,    282.05,  282.05,  282.05,
  281.9,     281.9,   281.9,   281.9,
  281.8,     281.8,   281.8,   281.8,
  281.75,    281.75,  281.75,  281.75,
  281.8,     281.8,   281.8,   281.8,
  281.9,     281.9,   281.9,   281.9,
  281.9,     281.9,   281.9,   281.9,
  281.45,    281.45,  281.45,  281.45,
  280.65,    280.65,  280.65,  280.65,
  280.2,     280.2,   280.2,   280.2,
  280.05,    280.05,  280.05,  280.05,
  279.7,     279.7,   279.7,   279.7,
  279.35,    279.35,  279.35,  279.35,
  279.15,    279.15,  279.15,  279.15,
  279,       279,     279,     279,
  278.9,     278.9,   278.9,   278.9,
  278.8,     278.8,   278.8,   278.8,
  278.65,    278.65,  278.65,  278.65,
  278.4,     278.4,   278.4,   278.4,
  277.95,    277.95,  277.95,  277.95,
  277.45,    277.45,  277.45,  277.45,
  276.85,    276.85,  276.85,  276.85,
  276.25,    276.25,  276.25,  276.25,
  275.85,    275.85,  275.85,  275.85,
  275.4,     275.4,   275.4,   275.4,
  274.85,    274.85,  274.85,  274.85,
  274.2,     274.2,   274.2,   274.2,
  273.6,     273.6,   273.6,   273.6,
  273.2,     273.2,   273.2,   273.2,
  273,       273,     273,     273,
  272.9,     272.9,   272.9,   272.9,
  272.9,     272.9,   272.9,   272.9,
  272.75,    272.75,  272.75,  272.75,
  272.4,     272.4,   272.4,   272.4,
  272.3,     272.3,   272.3,   272.3,
  272.25,    272.25,  272.25,  272.25,
  272.1,     272.1,   272.1,   272.1,
  272.1,     272.1,   272.1,   272.1,
  272.25,    272.25,  272.25,  272.25,
  272.5,     272.5,   272.5,   272.5,
  272.75,    272.75,  272.75,  272.75,
  272.85,    272.85,  272.85,  272.85,
  273.1,     273.1,   273.1,   273.1,
  273.95,    273.95,  273.95,  273.95,
  274.95,    274.95,  274.95,  274.95,
  276.1,     276.1,   276.1,   276.1,
  277.35,    277.35,  277.35,  277.35,
  278,       278,     278,     278,
  278.75,    278.75,  278.75,  278.75,
  279.45,    279.45,  279.45,  279.45,
  279.55,    279.55,  279.55,  279.55,
  279.1,     279.1,   279.1,   279.1,
  278.4,     278.4,   278.4,   278.4,
  277.9,     277.9,   277.9,   277.9,
  277.45,    277.45,  277.45,  277.45,
  276.95,    276.95,  276.95,  276.95,
  276.45,    276.45,  276.45,  276.45,
  276,       276,     276,     276,
  275.7,     275.7,   275.7,   275.7,
  275.65,    275.65,  275.65,  275.65,
  275.65,    275.65,  275.65,  275.65,
  275.5,     275.5,   275.5,   275.5,
  275.65,    275.65,  275.65,  275.65,
  276.3,     276.3,   276.3,   276.3,
  276.9,     276.9,   276.9,   276.9,
  277.35,    277.35,  277.35,  277.35,
  277.75,    277.75,  277.75,  277.75,
  278.1,     278.1,   278.1,   278.1,
  278.25,    278.25,  278.25,  278.25,
  278.3,     278.3,   278.3,   278.3,
  278.45,    278.45,  278.45,  278.45,
  278.7,     278.7,   278.7,   278.7,
  278.9,     278.9,   278.9,   278.9,
  279,       279,     279,     279,
  279.05,    279.05,  279.05,  279.05,
  279.05,    279.05,  279.05,  279.05,
  278.95,    278.95,  278.95,  278.95,
  278.85,    278.85,  278.85,  278.85,
  278.8,     278.8,   278.8,   278.8,
  278.7,     278.7,   278.7,   278.7,
  278.7,     278.7,   278.7,   278.7,
  278.65,    278.65,  278.65,  278.65,
  278.4,     278.4,   278.4,   278.4,
  278.05,    278.05,  278.05,  278.05,
  277.85,    277.85,  277.85,  277.85,
  278.1,     278.1,   278.1,   278.1,
  278.65,    278.65,  278.65,  278.65,
  279.45,    279.45,  279.45,  279.45,
  280.3,     280.3,   280.3,   280.3,
  280.9,     280.9,   280.9,   280.9,
  281.3,     281.3,   281.3,   281.3,
  281.45,    281.45,  281.45,  281.45,
  281.7,     281.7,   281.7,   281.7,
  282.15,    282.15,  282.15,  282.15,
  282.7,     282.7,   282.7,   282.7,
  283.15,    283.15,  283.15,  283.15,
  283.2,     283.2,   283.2,   283.2,
  283,       283,     283,     283,
  282.7,     282.7,   282.7,   282.7,
  282.55,    282.55,  282.55,  282.55,
  282.6,     282.6,   282.6,   282.6,
  282.65,    282.65,  282.65,  282.65,
  282.6,     282.6,   282.6,   282.6,
  282.4,     282.4,   282.4,   282.4,
  282.25,    282.25,  282.25,  282.25,
  282.15,    282.15,  282.15,  282.15,
  281.9,     281.9,   281.9,   281.9,
  281.7,     281.7,   281.7,   281.7,
  281.6,     281.6,   281.6,   281.6,
  281.6,     281.6,   281.6,   281.6,
  281.6,     281.6,   281.6,   281.6,
  281.5,     281.5,   281.5,   281.5,
  281.5,     281.5,   281.5,   281.5,
  281.5,     281.5,   281.5,   281.5,
  281.45,    281.45,  281.45,  281.45,
  281.55,    281.55,  281.55,  281.55,
  281.6,     281.6,   281.6,   281.6,
  281.45,    281.45,  281.45,  281.45,
  281.2,     281.2,   281.2,   281.2,
  280.95,    280.95,  280.95,  280.95,
  280.75,    280.75,  280.75,  280.75,
  280.6,     280.6,   280.6,   280.6,
  280.6,     280.6,   280.6,   280.6,
  280.55,    280.55,  280.55,  280.55,
  280.4,     280.4,   280.4,   280.4,
  280.15,    280.15,  280.15,  280.15,
  279.85,    279.85,  279.85,  279.85,
  279.7,     279.7,   279.7,   279.7,
  279.45,    279.45,  279.45,  279.45,
  279.15,    279.15,  279.15,  279.15,
  279.1,     279.1,   279.1,   279.1,
  279.25,    279.25,  279.25,  279.25,
  279.4,     279.4,   279.4,   279.4,
  279.55,    279.55,  279.55,  279.55,
  279.85,    279.85,  279.85,  279.85,
  280.2,     280.2,   280.2,   280.2,
  280.45,    280.45,  280.45,  280.45,
  280.7,     280.7,   280.7,   280.7,
  280.9,     280.9,   280.9,   280.9,
  281.1,     281.1,   281.1,   281.1,
  281.3,     281.3,   281.3,   281.3,
  281.45,    281.45,  281.45,  281.45,
  281.6,     281.6,   281.6,   281.6,
  281.65,    281.65,  281.65,  281.65,
  281.65,    281.65,  281.65,  281.65,
  281.6,     281.6,   281.6,   281.6,
  281.65,    281.65,  281.65,  281.65,
  281.6,     281.6,   281.6,   281.6,
  281.5,     281.5,   281.5,   281.5,
  281.6,     281.6,   281.6,   281.6,
  281.65,    281.65,  281.65,  281.65,
  281.7,     281.7,   281.7,   281.7,
  281.85,    281.85,  281.85,  281.85,
  282,       282,     282,     282,
  281.55,    281.55,  281.55,  281.55,
  280.8,     280.8,   280.8,   280.8,
  280.35,    280.35,  280.35,  280.35,
  279.9,     279.9,   279.9,   279.9,
  279.5,     279.5,   279.5,   279.5,
  279.25,    279.25,  279.25,  279.25,
  279,       279,     279,     279,
  278.7,     278.7,   278.7,   278.7,
  278.45,    278.45,  278.45,  278.45,
  278.3,     278.3,   278.3,   278.3,
  278.25,    278.25,  278.25,  278.25,
  278.2,     278.2,   278.2,   278.2,
  278,       278,     278,     278,
  277.85,    277.85,  277.85,  277.85,
  277.8,     277.8,   277.8,   277.8,
  277.6,     277.6,   277.6,   277.6,
  277.2,     277.2,   277.2,   277.2,
  276.7,     276.7,   276.7,   276.7,
  276.25,    276.25,  276.25,  276.25,
  276.05,    276.05,  276.05,  276.05,
  276.15,    276.15,  276.15,  276.15,
  276.3,     276.3,   276.3,   276.3,
  276.3,     276.3,   276.3,   276.3,
  276.1,     276.1,   276.1,   276.1,
  275.95,    275.95,  275.95,  275.95,
  276.05,    276.05,  276.05,  276.05,
  276.35,    276.35,  276.35,  276.35,
  276.9,     276.9,   276.9,   276.9,
  277.6,     277.6,   277.6,   277.6,
  278.1,     278.1,   278.1,   278.1,
  278.55,    278.55,  278.55,  278.55,
  279.2,     279.2,   279.2,   279.2,
  279.85,    279.85,  279.85,  279.85,
  280.1,     280.1,   280.1,   280.1,
  280.05,    280.05,  280.05,  280.05,
  280.25,    280.25,  280.25,  280.25,
  280.7,     280.7,   280.7,   280.7,
  280.95,    280.95,  280.95,  280.95,
  280.9,     280.9,   280.9,   280.9,
  280.75,    280.75,  280.75,  280.75,
  280.65,    280.65,  280.65,  280.65,
  280.6,     280.6,   280.6,   280.6,
  280.55,    280.55,  280.55,  280.55,
  280.5,     280.5,   280.5,   280.5,
  280.3,     280.3,   280.3,   280.3,
  280.05,    280.05,  280.05,  280.05,
  279.85,    279.85,  279.85,  279.85,
  279.6,     279.6,   279.6,   279.6,
  279.35,    279.35,  279.35,  279.35,
  279.25,    279.25,  279.25,  279.25,
  279.35,    279.35,  279.35,  279.35,
  279.5,     279.5,   279.5,   279.5,
  279.55,    279.55,  279.55,  279.55,
  279.35,    279.35,  279.35,  279.35,
  279.05,    279.05,  279.05,  279.05,
  278.7,     278.7,   278.7,   278.7,
  278.3,     278.3,   278.3,   278.3,
  278.1,     278.1,   278.1,   278.1,
  278.05,    278.05,  278.05,  278.05,
  278.15,    278.15,  278.15,  278.15,
  278.35,    278.35,  278.35,  278.35,
  278.55,    278.55,  278.55,  278.55,
  278.85,    278.85,  278.85,  278.85,
  279.35,    279.35,  279.35,  279.35,
  279.95,    279.95,  279.95,  279.95,
  280.65,    280.65,  280.65,  280.65,
  281.5,     281.5,   281.5,   281.5,
  282.25,    282.25,  282.25,  282.25,
  282.65,    282.65,  282.65,  282.65,
  282.7,     282.7,   282.7,   282.7,
  282.7,     282.7,   282.7,   282.7,
  282.55,    282.55,  282.55,  282.55,
  282.3,     282.3,   282.3,   282.3,
  282.25,    282.25,  282.25,  282.25,
  282.15,    282.15,  282.15,  282.15,
  282,       282,     282,     282,
  281.9,     281.9,   281.9,   281.9,
  281.9,     281.9,   281.9,   281.9,
  282.05,    282.05,  282.05,  282.05,
  282.15,    282.15,  282.15,  282.15,
  282.1,     282.1,   282.1,   282.1,
  282.05,    282.05,  282.05,  282.05,
  282.15,    282.15,  282.15,  282.15,
  282.4,     282.4,   282.4,   282.4,
  282.6,     282.6,   282.6,   282.6,
  282.75,    282.75,  282.75,  282.75,
  282.9,     282.9,   282.9,   282.9,
  283.15,    283.15,  283.15,  283.15,
  283.55,    283.55,  283.55,  283.55,
  283.85,    283.85,  283.85,  283.85,
  283.85,    283.85,  283.85,  283.85,
  283.55,    283.55,  283.55,  283.55,
  283.4,     283.4,   283.4,   283.4,
  283.4,     283.4,   283.4,   283.4,
  283.45,    283.45,  283.45,  283.45,
  283.25,    283.25,  283.25,  283.25,
  282.8,     282.8,   282.8,   282.8,
  282.65,    282.65,  282.65,  282.65,
  282.65,    282.65,  282.65,  282.65,
  282.65,    282.65,  282.65,  282.65,
  282.6,     282.6,   282.6,   282.6,
  282.55,    282.55,  282.55,  282.55,
  282.55,    282.55,  282.55,  282.55,
  282.6,     282.6,   282.6,   282.6,
  282.6,     282.6,   282.6,   282.6,
  282.55,    282.55,  282.55,  282.55,
  282.5,     282.5,   282.5,   282.5,
  282.45,    282.45,  282.45,  282.45,
  282.4,     282.4,   282.4,   282.4,
  282.35,    282.35,  282.35,  282.35,
  282.35,    282.35,  282.35,  282.35,
  282.3,     282.3,   282.3,   282.3,
  282,       282,     282,     282,
  281.65,    281.65,  281.65,  281.65,
  281.3,     281.3,   281.3,   281.3,
  280.9,     280.9,   280.9,   280.9,
  280.6,     280.6,   280.6,   280.6,
  280.3,     280.3,   280.3,   280.3,
  280,       280,     280,     280,
  279.8,     279.8,   279.8,   279.8,
  279.85,    279.85,  279.85,  279.85,
  279.85,    279.85,  279.85,  279.85,
  279.55,    279.55,  279.55,  279.55,
  279.35,    279.35,  279.35,  279.35,
  279.35,    279.35,  279.35,  279.35,
  279.4,     279.4,   279.4,   279.4,
  279.4,     279.4,   279.4,   279.4,
  279.45,    279.45,  279.45,  279.45,
  279.55,    279.55,  279.55,  279.55,
  279.4,     279.4,   279.4,   279.4,
  278.8,     278.8,   278.8,   278.8,
  278.6,     278.6,   278.6,   278.6,
  278.7,     278.7,   278.7,   278.7,
  278.1,     278.1,   278.1,   278.1,
  277.25,    277.25,  277.25,  277.25,
  276.95,    276.95,  276.95,  276.95,
  276.75,    276.75,  276.75,  276.75,
  276.95,    276.95,  276.95,  276.95,
  277.9,     277.9,   277.9,   277.9,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.4,     278.4,   278.4,   278.4,
  278.5,     278.5,   278.5,   278.5,
  278.6,     278.6,   278.6,   278.6,
  278.75,    278.75,  278.75,  278.75,
  278.9,     278.9,   278.9,   278.9,
  278.95,    278.95,  278.95,  278.95,
  279,       279,     279,     279,
  279.05,    279.05,  279.05,  279.05,
  279,       279,     279,     279,
  278.95,    278.95,  278.95,  278.95,
  278.9,     278.9,   278.9,   278.9,
  278.7,     278.7,   278.7,   278.7,
  278.55,    278.55,  278.55,  278.55,
  278.45,    278.45,  278.45,  278.45,
  278.3,     278.3,   278.3,   278.3,
  278.15,    278.15,  278.15,  278.15,
  277.9,     277.9,   277.9,   277.9,
  277.5,     277.5,   277.5,   277.5,
  277,       277,     277,     277,
  276.6,     276.6,   276.6,   276.6,
  276.3,     276.3,   276.3,   276.3,
  275.95,    275.95,  275.95,  275.95,
  275.65,    275.65,  275.65,  275.65,
  275.5,     275.5,   275.5,   275.5,
  275.3,     275.3,   275.3,   275.3,
  275.15,    275.15,  275.15,  275.15,
  275.05,    275.05,  275.05,  275.05,
  274.8,     274.8,   274.8,   274.8,
  274.6,     274.6,   274.6,   274.6,
  274.65,    274.65,  274.65,  274.65,
  275.05,    275.05,  275.05,  275.05,
  275.6,     275.6,   275.6,   275.6,
  276.2,     276.2,   276.2,   276.2,
  276.85,    276.85,  276.85,  276.85,
  277.3,     277.3,   277.3,   277.3,
  277.85,    277.85,  277.85,  277.85,
  278.6,     278.6,   278.6,   278.6,
  279.2,     279.2,   279.2,   279.2,
  279.35,    279.35,  279.35,  279.35,
  279.5,     279.5,   279.5,   279.5,
  279.65,    279.65,  279.65,  279.65,
  279.55,    279.55,  279.55,  279.55,
  279.55,    279.55,  279.55,  279.55,
  279.25,    279.25,  279.25,  279.25,
  279.15,    279.15,  279.15,  279.15,
  279.05,    279.05,  279.05,  279.05,
  278.3,     278.3,   278.3,   278.3,
  277.45,    277.45,  277.45,  277.45,
  276.75,    276.75,  276.75,  276.75,
  276.25,    276.25,  276.25,  276.25,
  276,       276,     276,     276,
  275.8,     275.8,   275.8,   275.8,
  275.35,    275.35,  275.35,  275.35,
  274.55,    274.55,  274.55,  274.55,
  273.75,    273.75,  273.75,  273.75,
  273.3,     273.3,   273.3,   273.3,
  273.5,     273.5,   273.5,   273.5,
  273.7,     273.7,   273.7,   273.7,
  273.3,     273.3,   273.3,   273.3,
  273.1,     273.1,   273.1,   273.1,
  273.15,    273.15,  273.15,  273.15,
  273.3,     273.3,   273.3,   273.3,
  273.55,    273.55,  273.55,  273.55,
  273.7,     273.7,   273.7,   273.7,
  273.85,    273.85,  273.85,  273.85,
  274,       274,     274,     274,
  273.95,    273.95,  273.95,  273.95,
  274.05,    274.05,  274.05,  274.05,
  274.4,     274.4,   274.4,   274.4,
  274.6,     274.6,   274.6,   274.6,
  274.75,    274.75,  274.75,  274.75,
  274.75,    274.75,  274.75,  274.75,
  274.6,     274.6,   274.6,   274.6,
  274.5,     274.5,   274.5,   274.5,
  274.4,     274.4,   274.4,   274.4,
  274.35,    274.35,  274.35,  274.35,
  274.4,     274.4,   274.4,   274.4,
  274.55,    274.55,  274.55,  274.55,
  274.8,     274.8,   274.8,   274.8,
  275.25,    275.25,  275.25,  275.25,
  276.1,     276.1,   276.1,   276.1,
  277.15,    277.15,  277.15,  277.15,
  278.05,    278.05,  278.05,  278.05,
  278.7,     278.7,   278.7,   278.7,
  279.25,    279.25,  279.25,  279.25,
  279.65,    279.65,  279.65,  279.65,
  279.75,    279.75,  279.75,  279.75,
  279.9,     279.9,   279.9,   279.9,
  280.05,    280.05,  280.05,  280.05,
  279.8,     279.8,   279.8,   279.8,
  279.9,     279.9,   279.9,   279.9,
  280.35,    280.35,  280.35,  280.35,
  280.2,     280.2,   280.2,   280.2,
  279.65,    279.65,  279.65,  279.65,
  279,       279,     279,     279,
  278.2,     278.2,   278.2,   278.2,
  277.4,     277.4,   277.4,   277.4,
  276.85,    276.85,  276.85,  276.85,
  276.65,    276.65,  276.65,  276.65,
  276.55,    276.55,  276.55,  276.55,
  276.2,     276.2,   276.2,   276.2,
  275.75,    275.75,  275.75,  275.75,
  275.6,     275.6,   275.6,   275.6,
  275.5,     275.5,   275.5,   275.5,
  275.2,     275.2,   275.2,   275.2,
  275.1,     275.1,   275.1,   275.1,
  275.3,     275.3,   275.3,   275.3,
  275.55,    275.55,  275.55,  275.55,
  275.7,     275.7,   275.7,   275.7,
  275.7,     275.7,   275.7,   275.7,
  275.6,     275.6,   275.6,   275.6,
  275.3,     275.3,   275.3,   275.3,
  274.9,     274.9,   274.9,   274.9,
  274.7,     274.7,   274.7,   274.7,
  274.4,     274.4,   274.4,   274.4,
  273.8,     273.8,   273.8,   273.8,
  273.45,    273.45,  273.45,  273.45,
  273.55,    273.55,  273.55,  273.55,
  273.65,    273.65,  273.65,  273.65,
  273.65,    273.65,  273.65,  273.65,
  273.7,     273.7,   273.7,   273.7,
  273.8,     273.8,   273.8,   273.8,
  273.85,    273.85,  273.85,  273.85,
  273.8,     273.8,   273.8,   273.8,
  273.75,    273.75,  273.75,  273.75,
  273.85,    273.85,  273.85,  273.85,
  274.2,     274.2,   274.2,   274.2,
  274.65,    274.65,  274.65,  274.65,
  275.15,    275.15,  275.15,  275.15,
  275.7,     275.7,   275.7,   275.7,
  276.25,    276.25,  276.25,  276.25,
  276.9,     276.9,   276.9,   276.9,
  277.5,     277.5,   277.5,   277.5,
  277.85,    277.85,  277.85,  277.85,
  278.1,     278.1,   278.1,   278.1,
  278.4,     278.4,   278.4,   278.4,
  278.65,    278.65,  278.65,  278.65,
  278.85,    278.85,  278.85,  278.85,
  278.85,    278.85,  278.85,  278.85,
  278.65,    278.65,  278.65,  278.65,
  278.5,     278.5,   278.5,   278.5,
  278.3,     278.3,   278.3,   278.3,
  277.95,    277.95,  277.95,  277.95,
  277.6,     277.6,   277.6,   277.6,
  277.3,     277.3,   277.3,   277.3,
  277.05,    277.05,  277.05,  277.05,
  276.95,    276.95,  276.95,  276.95,
  276.95,    276.95,  276.95,  276.95,
  276.85,    276.85,  276.85,  276.85,
  276.6,     276.6,   276.6,   276.6,
  276.35,    276.35,  276.35,  276.35,
  276.35,    276.35,  276.35,  276.35,
  276.6,     276.6,   276.6,   276.6,
  276.8,     276.8,   276.8,   276.8,
  276.8,     276.8,   276.8,   276.8,
  276.8,     276.8,   276.8,   276.8,
  276.85,    276.85,  276.85,  276.85,
  276.8,     276.8,   276.8,   276.8,
  276.8,     276.8,   276.8,   276.8,
  276.4,     276.4,   276.4,   276.4,
  275.45,    275.45,  275.45,  275.45,
  274.95,    274.95,  274.95,  274.95,
  275.1,     275.1,   275.1,   275.1,
  275.35,    275.35,  275.35,  275.35,
  275.6,     275.6,   275.6,   275.6,
  275.8,     275.8,   275.8,   275.8,
  275.95,    275.95,  275.95,  275.95,
  276.25,    276.25,  276.25,  276.25,
  276.55,    276.55,  276.55,  276.55,
  276.7,     276.7,   276.7,   276.7,
  276.7,     276.7,   276.7,   276.7,
  276.65,    276.65,  276.65,  276.65,
  276.7,     276.7,   276.7,   276.7,
  276.85,    276.85,  276.85,  276.85,
  277.05,    277.05,  277.05,  277.05,
  277.3,     277.3,   277.3,   277.3,
  277.7,     277.7,   277.7,   277.7,
  278.05,    278.05,  278.05,  278.05,
  278.3,     278.3,   278.3,   278.3,
  278.75,    278.75,  278.75,  278.75,
  279.2,     279.2,   279.2,   279.2,
  279.45,    279.45,  279.45,  279.45,
  279.85,    279.85,  279.85,  279.85,
  280.35,    280.35,  280.35,  280.35,
  280.7,     280.7,   280.7,   280.7,
  281.1,     281.1,   281.1,   281.1,
  281.45,    281.45,  281.45,  281.45,
  281.55,    281.55,  281.55,  281.55,
  281.6,     281.6,   281.6,   281.6,
  281.65,    281.65,  281.65,  281.65,
  281.65,    281.65,  281.65,  281.65,
  281.6,     281.6,   281.6,   281.6,
  281.5,     281.5,   281.5,   281.5,
  281.35,    281.35,  281.35,  281.35,
  281.2,     281.2,   281.2,   281.2,
  281.1,     281.1,   281.1,   281.1,
  281.1,     281.1,   281.1,   281.1,
  281.1,     281.1,   281.1,   281.1,
  281,       281,     281,     281,
  281,       281,     281,     281,
  281.15,    281.15,  281.15,  281.15,
  281.3,     281.3,   281.3,   281.3,
  281.35,    281.35,  281.35,  281.35,
  281.45,    281.45,  281.45,  281.45,
  281.4,     281.4,   281.4,   281.4,
  281,       281,     281,     281,
  280.65,    280.65,  280.65,  280.65,
  280.55,    280.55,  280.55,  280.55,
  280.55,    280.55,  280.55,  280.55,
  280.65,    280.65,  280.65,  280.65,
  280.75,    280.75,  280.75,  280.75,
  280.85,    280.85,  280.85,  280.85,
  281,       281,     281,     281,
  281.05,    281.05,  281.05,  281.05,
  281.05,    281.05,  281.05,  281.05,
  281.1,     281.1,   281.1,   281.1,
  281.2,     281.2,   281.2,   281.2,
  281.3,     281.3,   281.3,   281.3,
  281.4,     281.4,   281.4,   281.4,
  281.55,    281.55,  281.55,  281.55,
  281.8,     281.8,   281.8,   281.8,
  282,       282,     282,     282,
  282.05,    282.05,  282.05,  282.05,
  282.05,    282.05,  282.05,  282.05,
  282.3,     282.3,   282.3,   282.3,
  282.9,     282.9,   282.9,   282.9,
  283.15,    283.15,  283.15,  283.15,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283,       283,     283,     283,
  282.7,     282.7,   282.7,   282.7,
  282.25,    282.25,  282.25,  282.25,
  281.9,     281.9,   281.9,   281.9,
  281.8,     281.8,   281.8,   281.8,
  281.8,     281.8,   281.8,   281.8,
  281.75,    281.75,  281.75,  281.75,
  280.95,    280.95,  280.95,  280.95,
  279.35,    279.35,  279.35,  279.35,
  278.65,    278.65,  278.65,  278.65,
  278.65,    278.65,  278.65,  278.65,
  278.35,    278.35,  278.35,  278.35,
  277.95,    277.95,  277.95,  277.95,
  277.65,    277.65,  277.65,  277.65,
  277.55,    277.55,  277.55,  277.55,
  277.65,    277.65,  277.65,  277.65,
  278,       278,     278,     278,
  278.35,    278.35,  278.35,  278.35,
  278.5,     278.5,   278.5,   278.5,
  278.35,    278.35,  278.35,  278.35,
  278.2,     278.2,   278.2,   278.2,
  278.1,     278.1,   278.1,   278.1,
  277.85,    277.85,  277.85,  277.85,
  277.7,     277.7,   277.7,   277.7,
  277.6,     277.6,   277.6,   277.6,
  277.45,    277.45,  277.45,  277.45,
  277.45,    277.45,  277.45,  277.45,
  277.6,     277.6,   277.6,   277.6,
  277.55,    277.55,  277.55,  277.55,
  277.3,     277.3,   277.3,   277.3,
  277.1,     277.1,   277.1,   277.1,
  277,       277,     277,     277,
  276.95,    276.95,  276.95,  276.95,
  276.9,     276.9,   276.9,   276.9,
  276.65,    276.65,  276.65,  276.65,
  276.1,     276.1,   276.1,   276.1,
  275.5,     275.5,   275.5,   275.5,
  275,       275,     275,     275,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  275,       275,     275,     275,
  275.55,    275.55,  275.55,  275.55,
  276.3,     276.3,   276.3,   276.3,
  277.05,    277.05,  277.05,  277.05,
  277.55,    277.55,  277.55,  277.55,
  278.05,    278.05,  278.05,  278.05,
  278.55,    278.55,  278.55,  278.55,
  278.8,     278.8,   278.8,   278.8,
  278.9,     278.9,   278.9,   278.9,
  279,       279,     279,     279,
  279.1,     279.1,   279.1,   279.1,
  279.2,     279.2,   279.2,   279.2,
  279.25,    279.25,  279.25,  279.25,
  279.3,     279.3,   279.3,   279.3,
  279.4,     279.4,   279.4,   279.4,
  279.45,    279.45,  279.45,  279.45,
  279.45,    279.45,  279.45,  279.45,
  279.45,    279.45,  279.45,  279.45,
  279.5,     279.5,   279.5,   279.5,
  279.5,     279.5,   279.5,   279.5,
  279.4,     279.4,   279.4,   279.4,
  279.4,     279.4,   279.4,   279.4,
  279.5,     279.5,   279.5,   279.5,
  279.65,    279.65,  279.65,  279.65,
  279.7,     279.7,   279.7,   279.7,
  279.85,    279.85,  279.85,  279.85,
  279.85,    279.85,  279.85,  279.85,
  279.6,     279.6,   279.6,   279.6,
  279.55,    279.55,  279.55,  279.55,
  279.75,    279.75,  279.75,  279.75,
  280.25,    280.25,  280.25,  280.25,
  280.9,     280.9,   280.9,   280.9,
  281.3,     281.3,   281.3,   281.3,
  281.2,     281.2,   281.2,   281.2,
  281.1,     281.1,   281.1,   281.1,
  280.35,    280.35,  280.35,  280.35,
  279.1,     279.1,   279.1,   279.1,
  278.95,    278.95,  278.95,  278.95,
  279.3,     279.3,   279.3,   279.3,
  279.25,    279.25,  279.25,  279.25,
  279.15,    279.15,  279.15,  279.15,
  279.15,    279.15,  279.15,  279.15,
  279.15,    279.15,  279.15,  279.15,
  279.2,     279.2,   279.2,   279.2,
  279.25,    279.25,  279.25,  279.25,
  279.25,    279.25,  279.25,  279.25,
  279.2,     279.2,   279.2,   279.2,
  279.1,     279.1,   279.1,   279.1,
  279.15,    279.15,  279.15,  279.15,
  279.45,    279.45,  279.45,  279.45,
  279.85,    279.85,  279.85,  279.85,
  280.25,    280.25,  280.25,  280.25,
  280.65,    280.65,  280.65,  280.65,
  281.1,     281.1,   281.1,   281.1,
  281.4,     281.4,   281.4,   281.4,
  281.55,    281.55,  281.55,  281.55,
  281.65,    281.65,  281.65,  281.65,
  281.7,     281.7,   281.7,   281.7,
  281.8,     281.8,   281.8,   281.8,
  281.95,    281.95,  281.95,  281.95,
  282.1,     282.1,   282.1,   282.1,
  282.3,     282.3,   282.3,   282.3,
  282.55,    282.55,  282.55,  282.55,
  282.65,    282.65,  282.65,  282.65,
  282.55,    282.55,  282.55,  282.55,
  282.45,    282.45,  282.45,  282.45,
  282.4,     282.4,   282.4,   282.4,
  282.3,     282.3,   282.3,   282.3,
  282.3,     282.3,   282.3,   282.3,
  282.3,     282.3,   282.3,   282.3,
  282.2,     282.2,   282.2,   282.2,
  282.05,    282.05,  282.05,  282.05,
  281.95,    281.95,  281.95,  281.95,
  281.95,    281.95,  281.95,  281.95,
  281.95,    281.95,  281.95,  281.95,
  281.9,     281.9,   281.9,   281.9,
  281.8,     281.8,   281.8,   281.8,
  281.8,     281.8,   281.8,   281.8,
  281.8,     281.8,   281.8,   281.8,
  281.65,    281.65,  281.65,  281.65,
  281.6,     281.6,   281.6,   281.6,
  281.7,     281.7,   281.7,   281.7,
  281.75,    281.75,  281.75,  281.75,
  281.8,     281.8,   281.8,   281.8,
  281.8,     281.8,   281.8,   281.8,
  281.7,     281.7,   281.7,   281.7,
  281.7,     281.7,   281.7,   281.7,
  281.8,     281.8,   281.8,   281.8,
  281.9,     281.9,   281.9,   281.9,
  282,       282,     282,     282,
  282.05,    282.05,  282.05,  282.05,
  282.1,     282.1,   282.1,   282.1,
  282.15,    282.15,  282.15,  282.15,
  282.15,    282.15,  282.15,  282.15,
  282.2,     282.2,   282.2,   282.2,
  282.25,    282.25,  282.25,  282.25,
  282.3,     282.3,   282.3,   282.3,
  282.45,    282.45,  282.45,  282.45,
  282.6,     282.6,   282.6,   282.6,
  282.7,     282.7,   282.7,   282.7,
  282.8,     282.8,   282.8,   282.8,
  282.9,     282.9,   282.9,   282.9,
  282.6,     282.6,   282.6,   282.6,
  282.15,    282.15,  282.15,  282.15,
  282.05,    282.05,  282.05,  282.05,
  282.2,     282.2,   282.2,   282.2,
  282.5,     282.5,   282.5,   282.5,
  282.8,     282.8,   282.8,   282.8,
  283,       283,     283,     283,
  283.25,    283.25,  283.25,  283.25,
  283.5,     283.5,   283.5,   283.5,
  283.65,    283.65,  283.65,  283.65,
  283.7,     283.7,   283.7,   283.7,
  283.6,     283.6,   283.6,   283.6,
  283.4,     283.4,   283.4,   283.4,
  282.95,    282.95,  282.95,  282.95,
  282.3,     282.3,   282.3,   282.3,
  281.9,     281.9,   281.9,   281.9,
  281.85,    281.85,  281.85,  281.85,
  281.85,    281.85,  281.85,  281.85,
  281.8,     281.8,   281.8,   281.8,
  281.7,     281.7,   281.7,   281.7,
  281.55,    281.55,  281.55,  281.55,
  281.35,    281.35,  281.35,  281.35,
  281.05,    281.05,  281.05,  281.05,
  280.8,     280.8,   280.8,   280.8,
  280.65,    280.65,  280.65,  280.65,
  280.45,    280.45,  280.45,  280.45,
  280.3,     280.3,   280.3,   280.3,
  280.1,     280.1,   280.1,   280.1,
  279.75,    279.75,  279.75,  279.75,
  279.45,    279.45,  279.45,  279.45,
  279.35,    279.35,  279.35,  279.35,
  279.25,    279.25,  279.25,  279.25,
  279.2,     279.2,   279.2,   279.2,
  279.35,    279.35,  279.35,  279.35,
  279.6,     279.6,   279.6,   279.6,
  279.8,     279.8,   279.8,   279.8,
  280,       280,     280,     280,
  280.25,    280.25,  280.25,  280.25,
  280.4,     280.4,   280.4,   280.4,
  280.5,     280.5,   280.5,   280.5,
  280.5,     280.5,   280.5,   280.5,
  280.5,     280.5,   280.5,   280.5,
  280.65,    280.65,  280.65,  280.65,
  280.85,    280.85,  280.85,  280.85,
  281.05,    281.05,  281.05,  281.05,
  281.3,     281.3,   281.3,   281.3,
  281.6,     281.6,   281.6,   281.6,
  281.9,     281.9,   281.9,   281.9,
  282.25,    282.25,  282.25,  282.25,
  282.75,    282.75,  282.75,  282.75,
  283.1,     283.1,   283.1,   283.1,
  283.3,     283.3,   283.3,   283.3,
  283.6,     283.6,   283.6,   283.6,
  283.9,     283.9,   283.9,   283.9,
  284.15,    284.15,  284.15,  284.15,
  284.3,     284.3,   284.3,   284.3,
  284.3,     284.3,   284.3,   284.3,
  284.25,    284.25,  284.25,  284.25,
  284.15,    284.15,  284.15,  284.15,
  284,       284,     284,     284,
  283.85,    283.85,  283.85,  283.85,
  283.65,    283.65,  283.65,  283.65,
  283.45,    283.45,  283.45,  283.45,
  283.3,     283.3,   283.3,   283.3,
  283.2,     283.2,   283.2,   283.2,
  283.1,     283.1,   283.1,   283.1,
  283.2,     283.2,   283.2,   283.2,
  283.4,     283.4,   283.4,   283.4,
  283.4,     283.4,   283.4,   283.4,
  283.4,     283.4,   283.4,   283.4,
  283.45,    283.45,  283.45,  283.45,
  283.45,    283.45,  283.45,  283.45,
  283.45,    283.45,  283.45,  283.45,
  283.4,     283.4,   283.4,   283.4,
  283.25,    283.25,  283.25,  283.25,
  283.1,     283.1,   283.1,   283.1,
  282.9,     282.9,   282.9,   282.9,
  282.7,     282.7,   282.7,   282.7,
  282.45,    282.45,  282.45,  282.45,
  281.95,    281.95,  281.95,  281.95,
  281.45,    281.45,  281.45,  281.45,
  281.3,     281.3,   281.3,   281.3,
  281.35,    281.35,  281.35,  281.35,
  281.05,    281.05,  281.05,  281.05,
  280.5,     280.5,   280.5,   280.5,
  280.15,    280.15,  280.15,  280.15,
  280,       280,     280,     280,
  279.95,    279.95,  279.95,  279.95,
  280.05,    280.05,  280.05,  280.05,
  280.4,     280.4,   280.4,   280.4,
  280.7,     280.7,   280.7,   280.7,
  280.85,    280.85,  280.85,  280.85,
  280.95,    280.95,  280.95,  280.95,
  281.15,    281.15,  281.15,  281.15,
  281.5,     281.5,   281.5,   281.5,
  281.95,    281.95,  281.95,  281.95,
  282.7,     282.7,   282.7,   282.7,
  283.4,     283.4,   283.4,   283.4,
  283.85,    283.85,  283.85,  283.85,
  284.1,     284.1,   284.1,   284.1,
  284.2,     284.2,   284.2,   284.2,
  284.45,    284.45,  284.45,  284.45,
  284.7,     284.7,   284.7,   284.7,
  284.75,    284.75,  284.75,  284.75,
  284.7,     284.7,   284.7,   284.7,
  284.65,    284.65,  284.65,  284.65,
  284.6,     284.6,   284.6,   284.6,
  284.55,    284.55,  284.55,  284.55,
  284.55,    284.55,  284.55,  284.55,
  284.55,    284.55,  284.55,  284.55,
  284.5,     284.5,   284.5,   284.5,
  284.35,    284.35,  284.35,  284.35,
  284.15,    284.15,  284.15,  284.15,
  283.85,    283.85,  283.85,  283.85,
  283.55,    283.55,  283.55,  283.55,
  283.35,    283.35,  283.35,  283.35,
  283.2,     283.2,   283.2,   283.2,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  283.2,     283.2,   283.2,   283.2,
  283.3,     283.3,   283.3,   283.3,
  283.3,     283.3,   283.3,   283.3,
  283.25,    283.25,  283.25,  283.25,
  283.3,     283.3,   283.3,   283.3,
  283.4,     283.4,   283.4,   283.4,
  283.4,     283.4,   283.4,   283.4,
  283.35,    283.35,  283.35,  283.35,
  283.3,     283.3,   283.3,   283.3,
  283.3,     283.3,   283.3,   283.3,
  283.45,    283.45,  283.45,  283.45,
  283.7,     283.7,   283.7,   283.7,
  283.9,     283.9,   283.9,   283.9,
  283.85,    283.85,  283.85,  283.85,
  283.25,    283.25,  283.25,  283.25,
  282.7,     282.7,   282.7,   282.7,
  282.75,    282.75,  282.75,  282.75,
  282.95,    282.95,  282.95,  282.95,
  283,       283,     283,     283,
  281.7,     281.7,   281.7,   281.7,
  280.75,    280.75,  280.75,  280.75,
  281.55,    281.55,  281.55,  281.55,
  282.2,     282.2,   282.2,   282.2,
  282.2,     282.2,   282.2,   282.2,
  281.9,     281.9,   281.9,   281.9,
  282.1,     282.1,   282.1,   282.1,
  282.6,     282.6,   282.6,   282.6,
  282.7,     282.7,   282.7,   282.7,
  282.5,     282.5,   282.5,   282.5,
  282.1,     282.1,   282.1,   282.1,
  281.4,     281.4,   281.4,   281.4,
  280.55,    280.55,  280.55,  280.55,
  280.05,    280.05,  280.05,  280.05,
  280.2,     280.2,   280.2,   280.2,
  280.8,     280.8,   280.8,   280.8,
  281.3,     281.3,   281.3,   281.3,
  281.3,     281.3,   281.3,   281.3,
  281.1,     281.1,   281.1,   281.1,
  281.1,     281.1,   281.1,   281.1,
  281.2,     281.2,   281.2,   281.2,
  281.25,    281.25,  281.25,  281.25,
  281.4,     281.4,   281.4,   281.4,
  281.45,    281.45,  281.45,  281.45,
  281.05,    281.05,  281.05,  281.05,
  280.8,     280.8,   280.8,   280.8,
  281,       281,     281,     281,
  281.75,    281.75,  281.75,  281.75,
  282.7,     282.7,   282.7,   282.7,
  283.25,    283.25,  283.25,  283.25,
  283.65,    283.65,  283.65,  283.65,
  284,       284,     284,     284,
  284.4,     284.4,   284.4,   284.4,
  284.8,     284.8,   284.8,   284.8,
  284.8,     284.8,   284.8,   284.8,
  284.95,    284.95,  284.95,  284.95,
  285.25,    285.25,  285.25,  285.25,
  285.15,    285.15,  285.15,  285.15,
  285,       285,     285,     285,
  284.75,    284.75,  284.75,  284.75,
  283.3,     283.3,   283.3,   283.3,
  282.35,    282.35,  282.35,  282.35,
  283.15,    283.15,  283.15,  283.15,
  283.7,     283.7,   283.7,   283.7,
  283.05,    283.05,  283.05,  283.05,
  281.95,    281.95,  281.95,  281.95,
  281.85,    281.85,  281.85,  281.85,
  282.65,    282.65,  282.65,  282.65,
  283.3,     283.3,   283.3,   283.3,
  283.25,    283.25,  283.25,  283.25,
  282.35,    282.35,  282.35,  282.35,
  282.2,     282.2,   282.2,   282.2,
  283.25,    283.25,  283.25,  283.25,
  284.2,     284.2,   284.2,   284.2,
  284.65,    284.65,  284.65,  284.65,
  284.55,    284.55,  284.55,  284.55,
  284.4,     284.4,   284.4,   284.4,
  284.4,     284.4,   284.4,   284.4,
  284.35,    284.35,  284.35,  284.35,
  284.15,    284.15,  284.15,  284.15,
  284.05,    284.05,  284.05,  284.05,
  283.95,    283.95,  283.95,  283.95,
  283.85,    283.85,  283.85,  283.85,
  283.9,     283.9,   283.9,   283.9,
  283.95,    283.95,  283.95,  283.95,
  283.85,    283.85,  283.85,  283.85,
  283.75,    283.75,  283.75,  283.75,
  283.7,     283.7,   283.7,   283.7,
  283.55,    283.55,  283.55,  283.55,
  283.3,     283.3,   283.3,   283.3,
  283.05,    283.05,  283.05,  283.05,
  282.95,    282.95,  282.95,  282.95,
  283,       283,     283,     283,
  283,       283,     283,     283,
  282.6,     282.6,   282.6,   282.6,
  282.1,     282.1,   282.1,   282.1,
  281.85,    281.85,  281.85,  281.85,
  281.55,    281.55,  281.55,  281.55,
  281.4,     281.4,   281.4,   281.4,
  281.6,     281.6,   281.6,   281.6,
  281.8,     281.8,   281.8,   281.8,
  281.9,     281.9,   281.9,   281.9,
  282.05,    282.05,  282.05,  282.05,
  282.15,    282.15,  282.15,  282.15,
  282.1,     282.1,   282.1,   282.1,
  282,       282,     282,     282,
  281.7,     281.7,   281.7,   281.7,
  281.45,    281.45,  281.45,  281.45,
  281.2,     281.2,   281.2,   281.2,
  280.75,    280.75,  280.75,  280.75,
  280.35,    280.35,  280.35,  280.35,
  280,       280,     280,     280,
  279.8,     279.8,   279.8,   279.8,
  279.85,    279.85,  279.85,  279.85,
  280.1,     280.1,   280.1,   280.1,
  280.45,    280.45,  280.45,  280.45,
  280.8,     280.8,   280.8,   280.8,
  280.65,    280.65,  280.65,  280.65,
  279.95,    279.95,  279.95,  279.95,
  279.75,    279.75,  279.75,  279.75,
  280,       280,     280,     280,
  279.8,     279.8,   279.8,   279.8,
  280.1,     280.1,   280.1,   280.1,
  280.65,    280.65,  280.65,  280.65,
  280.15,    280.15,  280.15,  280.15,
  279.5,     279.5,   279.5,   279.5,
  280.05,    280.05,  280.05,  280.05,
  281.05,    281.05,  281.05,  281.05,
  281.05,    281.05,  281.05,  281.05,
  280.8,     280.8,   280.8,   280.8,
  280.2,     280.2,   280.2,   280.2,
  279.95,    279.95,  279.95,  279.95,
  280.6,     280.6,   280.6,   280.6,
  280.25,    280.25,  280.25,  280.25,
  279.5,     279.5,   279.5,   279.5,
  279.4,     279.4,   279.4,   279.4,
  279.6,     279.6,   279.6,   279.6,
  279.75,    279.75,  279.75,  279.75,
  279.5,     279.5,   279.5,   279.5,
  279.05,    279.05,  279.05,  279.05,
  278.7,     278.7,   278.7,   278.7,
  278.55,    278.55,  278.55,  278.55,
  278.65,    278.65,  278.65,  278.65,
  278.85,    278.85,  278.85,  278.85,
  278.95,    278.95,  278.95,  278.95,
  278.95,    278.95,  278.95,  278.95,
  278.95,    278.95,  278.95,  278.95,
  278.9,     278.9,   278.9,   278.9,
  278.85,    278.85,  278.85,  278.85,
  278.85,    278.85,  278.85,  278.85,
  278.75,    278.75,  278.75,  278.75,
  278.4,     278.4,   278.4,   278.4,
  277.95,    277.95,  277.95,  277.95,
  277.5,     277.5,   277.5,   277.5,
  276.95,    276.95,  276.95,  276.95,
  276.45,    276.45,  276.45,  276.45,
  276.3,     276.3,   276.3,   276.3,
  276.25,    276.25,  276.25,  276.25,
  276,       276,     276,     276,
  275.75,    275.75,  275.75,  275.75,
  275.55,    275.55,  275.55,  275.55,
  275.4,     275.4,   275.4,   275.4,
  275.4,     275.4,   275.4,   275.4,
  275.65,    275.65,  275.65,  275.65,
  276.35,    276.35,  276.35,  276.35,
  277.4,     277.4,   277.4,   277.4,
  277.9,     277.9,   277.9,   277.9,
  277.9,     277.9,   277.9,   277.9,
  278.25,    278.25,  278.25,  278.25,
  278.9,     278.9,   278.9,   278.9,
  279.55,    279.55,  279.55,  279.55,
  280.05,    280.05,  280.05,  280.05,
  280.45,    280.45,  280.45,  280.45,
  280.75,    280.75,  280.75,  280.75,
  281,       281,     281,     281,
  281.15,    281.15,  281.15,  281.15,
  281.25,    281.25,  281.25,  281.25,
  281.4,     281.4,   281.4,   281.4,
  281.35,    281.35,  281.35,  281.35,
  281.05,    281.05,  281.05,  281.05,
  280.8,     280.8,   280.8,   280.8,
  280.6,     280.6,   280.6,   280.6,
  280.3,     280.3,   280.3,   280.3,
  280.1,     280.1,   280.1,   280.1,
  280.05,    280.05,  280.05,  280.05,
  280.05,    280.05,  280.05,  280.05,
  279.95,    279.95,  279.95,  279.95,
  279.85,    279.85,  279.85,  279.85,
  279.9,     279.9,   279.9,   279.9,
  280.2,     280.2,   280.2,   280.2,
  280.6,     280.6,   280.6,   280.6,
  280.7,     280.7,   280.7,   280.7,
  280.55,    280.55,  280.55,  280.55,
  280.35,    280.35,  280.35,  280.35,
  280.25,    280.25,  280.25,  280.25,
  280.25,    280.25,  280.25,  280.25,
  280.15,    280.15,  280.15,  280.15,
  280,       280,     280,     280,
  279.9,     279.9,   279.9,   279.9,
  279.85,    279.85,  279.85,  279.85,
  279.9,     279.9,   279.9,   279.9,
  279.95,    279.95,  279.95,  279.95,
  279.9,     279.9,   279.9,   279.9,
  279.8,     279.8,   279.8,   279.8,
  279.7,     279.7,   279.7,   279.7,
  279.6,     279.6,   279.6,   279.6,
  279.5,     279.5,   279.5,   279.5,
  279.45,    279.45,  279.45,  279.45,
  279.4,     279.4,   279.4,   279.4,
  279.35,    279.35,  279.35,  279.35,
  279.4,     279.4,   279.4,   279.4,
  279.65,    279.65,  279.65,  279.65,
  280.2,     280.2,   280.2,   280.2,
  280.95,    280.95,  280.95,  280.95,
  281.65,    281.65,  281.65,  281.65,
  282.3,     282.3,   282.3,   282.3,
  282.65,    282.65,  282.65,  282.65,
  282.8,     282.8,   282.8,   282.8,
  283.55,    283.55,  283.55,  283.55,
  284.35,    284.35,  284.35,  284.35,
  284.9,     284.9,   284.9,   284.9,
  285.6,     285.6,   285.6,   285.6,
  286.15,    286.15,  286.15,  286.15,
  286.45,    286.45,  286.45,  286.45,
  286.65,    286.65,  286.65,  286.65,
  286.9,     286.9,   286.9,   286.9,
  287,       287,     287,     287,
  286.85,    286.85,  286.85,  286.85,
  286.6,     286.6,   286.6,   286.6,
  286.25,    286.25,  286.25,  286.25,
  285.75,    285.75,  285.75,  285.75,
  285.2,     285.2,   285.2,   285.2,
  284.9,     284.9,   284.9,   284.9,
  284.75,    284.75,  284.75,  284.75,
  284.55,    284.55,  284.55,  284.55,
  284.35,    284.35,  284.35,  284.35,
  284.1,     284.1,   284.1,   284.1,
  283.6,     283.6,   283.6,   283.6,
  283.2,     283.2,   283.2,   283.2,
  283,       283,     283,     283,
  282.6,     282.6,   282.6,   282.6,
  282,       282,     282,     282,
  281.65,    281.65,  281.65,  281.65,
  281.7,     281.7,   281.7,   281.7,
  281.75,    281.75,  281.75,  281.75,
  281.75,    281.75,  281.75,  281.75,
  281.75,    281.75,  281.75,  281.75,
  281.7,     281.7,   281.7,   281.7,
  281.5,     281.5,   281.5,   281.5,
  281.1,     281.1,   281.1,   281.1,
  280.55,    280.55,  280.55,  280.55,
  279.95,    279.95,  279.95,  279.95,
  279.35,    279.35,  279.35,  279.35,
  278.8,     278.8,   278.8,   278.8,
  278.4,     278.4,   278.4,   278.4,
  278.05,    278.05,  278.05,  278.05,
  277.7,     277.7,   277.7,   277.7,
  277.45,    277.45,  277.45,  277.45,
  277.5,     277.5,   277.5,   277.5,
  277.95,    277.95,  277.95,  277.95,
  278.55,    278.55,  278.55,  278.55,
  279.35,    279.35,  279.35,  279.35,
  280.3,     280.3,   280.3,   280.3,
  281.2,     281.2,   281.2,   281.2,
  282.1,     282.1,   282.1,   282.1,
  282.9,     282.9,   282.9,   282.9,
  283.45,    283.45,  283.45,  283.45,
  283.85,    283.85,  283.85,  283.85,
  284.25,    284.25,  284.25,  284.25,
  284.55,    284.55,  284.55,  284.55,
  284.8,     284.8,   284.8,   284.8,
  285.1,     285.1,   285.1,   285.1,
  285.3,     285.3,   285.3,   285.3,
  285.45,    285.45,  285.45,  285.45,
  285.3,     285.3,   285.3,   285.3,
  285,       285,     285,     285,
  284.8,     284.8,   284.8,   284.8,
  284.5,     284.5,   284.5,   284.5,
  284.35,    284.35,  284.35,  284.35,
  284.35,    284.35,  284.35,  284.35,
  284.35,    284.35,  284.35,  284.35,
  284.35,    284.35,  284.35,  284.35,
  284.45,    284.45,  284.45,  284.45,
  284.65,    284.65,  284.65,  284.65,
  284.85,    284.85,  284.85,  284.85,
  285,       285,     285,     285,
  285,       285,     285,     285,
  284.9,     284.9,   284.9,   284.9,
  284.85,    284.85,  284.85,  284.85,
  284.8,     284.8,   284.8,   284.8,
  284.7,     284.7,   284.7,   284.7,
  284.7,     284.7,   284.7,   284.7,
  284.7,     284.7,   284.7,   284.7,
  284.65,    284.65,  284.65,  284.65,
  284.65,    284.65,  284.65,  284.65,
  284.6,     284.6,   284.6,   284.6,
  284.6,     284.6,   284.6,   284.6,
  284.75,    284.75,  284.75,  284.75,
  284.8,     284.8,   284.8,   284.8,
  284.7,     284.7,   284.7,   284.7,
  284.6,     284.6,   284.6,   284.6,
  284.45,    284.45,  284.45,  284.45,
  284.25,    284.25,  284.25,  284.25,
  284.05,    284.05,  284.05,  284.05,
  283.95,    283.95,  283.95,  283.95,
  283.95,    283.95,  283.95,  283.95,
  283.95,    283.95,  283.95,  283.95,
  283.95,    283.95,  283.95,  283.95,
  284,       284,     284,     284,
  284.1,     284.1,   284.1,   284.1,
  284.2,     284.2,   284.2,   284.2,
  284.3,     284.3,   284.3,   284.3,
  284.65,    284.65,  284.65,  284.65,
  285.15,    285.15,  285.15,  285.15,
  285.35,    285.35,  285.35,  285.35,
  285.2,     285.2,   285.2,   285.2,
  284.85,    284.85,  284.85,  284.85,
  284.35,    284.35,  284.35,  284.35,
  284,       284,     284,     284,
  284.1,     284.1,   284.1,   284.1,
  284.05,    284.05,  284.05,  284.05,
  283.3,     283.3,   283.3,   283.3,
  282.5,     282.5,   282.5,   282.5,
  282.15,    282.15,  282.15,  282.15,
  282.05,    282.05,  282.05,  282.05,
  282.05,    282.05,  282.05,  282.05,
  281.95,    281.95,  281.95,  281.95,
  281.5,     281.5,   281.5,   281.5,
  280.85,    280.85,  280.85,  280.85,
  280.55,    280.55,  280.55,  280.55,
  280.4,     280.4,   280.4,   280.4,
  280.1,     280.1,   280.1,   280.1,
  279.8,     279.8,   279.8,   279.8,
  279.6,     279.6,   279.6,   279.6,
  279.75,    279.75,  279.75,  279.75,
  279.95,    279.95,  279.95,  279.95,
  279.85,    279.85,  279.85,  279.85,
  279.7,     279.7,   279.7,   279.7,
  279.6,     279.6,   279.6,   279.6,
  279.5,     279.5,   279.5,   279.5,
  279.45,    279.45,  279.45,  279.45,
  279.4,     279.4,   279.4,   279.4,
  279.3,     279.3,   279.3,   279.3,
  279.2,     279.2,   279.2,   279.2,
  278.95,    278.95,  278.95,  278.95,
  278.55,    278.55,  278.55,  278.55,
  278.2,     278.2,   278.2,   278.2,
  277.95,    277.95,  277.95,  277.95,
  277.6,     277.6,   277.6,   277.6,
  277.3,     277.3,   277.3,   277.3,
  277.1,     277.1,   277.1,   277.1,
  276.9,     276.9,   276.9,   276.9,
  276.9,     276.9,   276.9,   276.9,
  276.85,    276.85,  276.85,  276.85,
  276.8,     276.8,   276.8,   276.8,
  277.05,    277.05,  277.05,  277.05,
  277.75,    277.75,  277.75,  277.75,
  278.5,     278.5,   278.5,   278.5,
  279.1,     279.1,   279.1,   279.1,
  279.85,    279.85,  279.85,  279.85,
  280.6,     280.6,   280.6,   280.6,
  281.25,    281.25,  281.25,  281.25,
  281.8,     281.8,   281.8,   281.8,
  282.2,     282.2,   282.2,   282.2,
  282.65,    282.65,  282.65,  282.65,
  282.9,     282.9,   282.9,   282.9,
  283,       283,     283,     283,
  283.15,    283.15,  283.15,  283.15,
  283,       283,     283,     283,
  282.75,    282.75,  282.75,  282.75,
  282.6,     282.6,   282.6,   282.6,
  282.45,    282.45,  282.45,  282.45,
  282.2,     282.2,   282.2,   282.2,
  281.9,     281.9,   281.9,   281.9,
  281.5,     281.5,   281.5,   281.5,
  281.15,    281.15,  281.15,  281.15,
  280.95,    280.95,  280.95,  280.95,
  280.55,    280.55,  280.55,  280.55,
  280.1,     280.1,   280.1,   280.1,
  279.75,    279.75,  279.75,  279.75,
  279.45,    279.45,  279.45,  279.45,
  279.1,     279.1,   279.1,   279.1,
  278.6,     278.6,   278.6,   278.6,
  278.5,     278.5,   278.5,   278.5,
  278.45,    278.45,  278.45,  278.45,
  278.3,     278.3,   278.3,   278.3,
  278.2,     278.2,   278.2,   278.2,
  277.85,    277.85,  277.85,  277.85,
  277.75,    277.75,  277.75,  277.75,
  277.85,    277.85,  277.85,  277.85,
  277.65,    277.65,  277.65,  277.65,
  277.45,    277.45,  277.45,  277.45,
  277.45,    277.45,  277.45,  277.45,
  277.45,    277.45,  277.45,  277.45,
  277.25,    277.25,  277.25,  277.25,
  276.85,    276.85,  276.85,  276.85,
  276.5,     276.5,   276.5,   276.5,
  276.2,     276.2,   276.2,   276.2,
  275.9,     275.9,   275.9,   275.9,
  275.6,     275.6,   275.6,   275.6,
  275.5,     275.5,   275.5,   275.5,
  275.55,    275.55,  275.55,  275.55,
  275.8,     275.8,   275.8,   275.8,
  276.6,     276.6,   276.6,   276.6,
  278,       278,     278,     278,
  279.35,    279.35,  279.35,  279.35,
  280.25,    280.25,  280.25,  280.25,
  280.95,    280.95,  280.95,  280.95,
  281.55,    281.55,  281.55,  281.55,
  282.05,    282.05,  282.05,  282.05,
  282.45,    282.45,  282.45,  282.45,
  282.8,     282.8,   282.8,   282.8,
  283.05,    283.05,  283.05,  283.05,
  283.4,     283.4,   283.4,   283.4,
  283.8,     283.8,   283.8,   283.8,
  284.05,    284.05,  284.05,  284.05,
  284.15,    284.15,  284.15,  284.15,
  284.3,     284.3,   284.3,   284.3,
  284.65,    284.65,  284.65,  284.65,
  284.7,     284.7,   284.7,   284.7,
  284.55,    284.55,  284.55,  284.55,
  284.4,     284.4,   284.4,   284.4,
  284.05,    284.05,  284.05,  284.05,
  283.75,    283.75,  283.75,  283.75,
  283.45,    283.45,  283.45,  283.45,
  283.15,    283.15,  283.15,  283.15,
  283.1,     283.1,   283.1,   283.1,
  283.15,    283.15,  283.15,  283.15,
  283.1,     283.1,   283.1,   283.1,
  282.95,    282.95,  282.95,  282.95,
  282.8,     282.8,   282.8,   282.8,
  282.65,    282.65,  282.65,  282.65,
  282.4,     282.4,   282.4,   282.4,
  282.2,     282.2,   282.2,   282.2,
  282.05,    282.05,  282.05,  282.05,
  281.95,    281.95,  281.95,  281.95,
  281.8,     281.8,   281.8,   281.8,
  281.5,     281.5,   281.5,   281.5,
  281.2,     281.2,   281.2,   281.2,
  281,       281,     281,     281,
  280.85,    280.85,  280.85,  280.85,
  280.65,    280.65,  280.65,  280.65,
  280.55,    280.55,  280.55,  280.55,
  280.55,    280.55,  280.55,  280.55,
  280.5,     280.5,   280.5,   280.5,
  280.45,    280.45,  280.45,  280.45,
  280.5,     280.5,   280.5,   280.5,
  280.6,     280.6,   280.6,   280.6,
  280.7,     280.7,   280.7,   280.7,
  280.9,     280.9,   280.9,   280.9,
  281.25,    281.25,  281.25,  281.25,
  281.65,    281.65,  281.65,  281.65,
  282.05,    282.05,  282.05,  282.05,
  282.35,    282.35,  282.35,  282.35,
  282.7,     282.7,   282.7,   282.7,
  283.25,    283.25,  283.25,  283.25,
  283.6,     283.6,   283.6,   283.6,
  283.15,    283.15,  283.15,  283.15,
  282.85,    282.85,  282.85,  282.85,
  283.25,    283.25,  283.25,  283.25,
  283.35,    283.35,  283.35,  283.35,
  283.15,    283.15,  283.15,  283.15,
  283.3,     283.3,   283.3,   283.3,
  283.75,    283.75,  283.75,  283.75,
  284,       284,     284,     284,
  284,       284,     284,     284,
  284,       284,     284,     284,
  283.95,    283.95,  283.95,  283.95,
  283.75,    283.75,  283.75,  283.75,
  283.4,     283.4,   283.4,   283.4,
  282.85,    282.85,  282.85,  282.85,
  282.2,     282.2,   282.2,   282.2,
  281.75,    281.75,  281.75,  281.75,
  281.75,    281.75,  281.75,  281.75,
  282,       282,     282,     282,
  282.05,    282.05,  282.05,  282.05,
  281.9,     281.9,   281.9,   281.9,
  281.7,     281.7,   281.7,   281.7,
  281.35,    281.35,  281.35,  281.35,
  280.8,     280.8,   280.8,   280.8,
  280.1,     280.1,   280.1,   280.1,
  279.6,     279.6,   279.6,   279.6,
  279.3,     279.3,   279.3,   279.3,
  279.25,    279.25,  279.25,  279.25,
  279.55,    279.55,  279.55,  279.55,
  279.85,    279.85,  279.85,  279.85,
  280.05,    280.05,  280.05,  280.05,
  280.25,    280.25,  280.25,  280.25,
  280.4,     280.4,   280.4,   280.4,
  280.4,     280.4,   280.4,   280.4,
  280.1,     280.1,   280.1,   280.1,
  279.65,    279.65,  279.65,  279.65,
  279.45,    279.45,  279.45,  279.45,
  279.45,    279.45,  279.45,  279.45,
  279.5,     279.5,   279.5,   279.5,
  279.6,     279.6,   279.6,   279.6,
  279.7,     279.7,   279.7,   279.7,
  279.85,    279.85,  279.85,  279.85,
  279.9,     279.9,   279.9,   279.9,
  279.8,     279.8,   279.8,   279.8,
  279.65,    279.65,  279.65,  279.65,
  279.55,    279.55,  279.55,  279.55,
  279.85,    279.85,  279.85,  279.85,
  280.5,     280.5,   280.5,   280.5,
  281,       281,     281,     281,
  281.6,     281.6,   281.6,   281.6,
  282.4,     282.4,   282.4,   282.4,
  283.1,     283.1,   283.1,   283.1,
  283.5,     283.5,   283.5,   283.5,
  283.45,    283.45,  283.45,  283.45,
  283.3,     283.3,   283.3,   283.3,
  283.4,     283.4,   283.4,   283.4,
  283.6,     283.6,   283.6,   283.6,
  283.55,    283.55,  283.55,  283.55,
  283.4,     283.4,   283.4,   283.4,
  283.1,     283.1,   283.1,   283.1,
  282.75,    282.75,  282.75,  282.75,
  282.65,    282.65,  282.65,  282.65,
  282.35,    282.35,  282.35,  282.35,
  281.7,     281.7,   281.7,   281.7,
  281.05,    281.05,  281.05,  281.05,
  280.3,     280.3,   280.3,   280.3,
  279.65,    279.65,  279.65,  279.65,
  279.1,     279.1,   279.1,   279.1,
  278.7,     278.7,   278.7,   278.7,
  278.5,     278.5,   278.5,   278.5,
  278.15,    278.15,  278.15,  278.15,
  277.9,     277.9,   277.9,   277.9,
  277.75,    277.75,  277.75,  277.75,
  277.6,     277.6,   277.6,   277.6,
  277.45,    277.45,  277.45,  277.45,
  277.3,     277.3,   277.3,   277.3,
  277.2,     277.2,   277.2,   277.2,
  277.15,    277.15,  277.15,  277.15,
  277.1,     277.1,   277.1,   277.1,
  276.95,    276.95,  276.95,  276.95,
  276.85,    276.85,  276.85,  276.85,
  276.7,     276.7,   276.7,   276.7,
  276.4,     276.4,   276.4,   276.4,
  276.3,     276.3,   276.3,   276.3,
  276.45,    276.45,  276.45,  276.45,
  276.7,     276.7,   276.7,   276.7,
  277.05,    277.05,  277.05,  277.05,
  277.35,    277.35,  277.35,  277.35,
  277.6,     277.6,   277.6,   277.6,
  277.9,     277.9,   277.9,   277.9,
  278.25,    278.25,  278.25,  278.25,
  278.65,    278.65,  278.65,  278.65,
  279.25,    279.25,  279.25,  279.25,
  280.25,    280.25,  280.25,  280.25,
  281.2,     281.2,   281.2,   281.2,
  281.9,     281.9,   281.9,   281.9,
  282.55,    282.55,  282.55,  282.55,
  283.35,    283.35,  283.35,  283.35,
  284.45,    284.45,  284.45,  284.45,
  285.45,    285.45,  285.45,  285.45,
  286,       286,     286,     286,
  286.35,    286.35,  286.35,  286.35,
  286.5,     286.5,   286.5,   286.5,
  286.5,     286.5,   286.5,   286.5,
  286.65,    286.65,  286.65,  286.65,
  286.95,    286.95,  286.95,  286.95,
  287.2,     287.2,   287.2,   287.2,
  287,       287,     287,     287,
  286.65,    286.65,  286.65,  286.65,
  286.4,     286.4,   286.4,   286.4,
  286,       286,     286,     286,
  285.55,    285.55,  285.55,  285.55,
  285.15,    285.15,  285.15,  285.15,
  284.7,     284.7,   284.7,   284.7,
  284.1,     284.1,   284.1,   284.1,
  283.5,     283.5,   283.5,   283.5,
  283,       283,     283,     283,
  282.5,     282.5,   282.5,   282.5,
  282.1,     282.1,   282.1,   282.1,
  281.8,     281.8,   281.8,   281.8,
  281.6,     281.6,   281.6,   281.6,
  281.5,     281.5,   281.5,   281.5,
  281.45,    281.45,  281.45,  281.45,
  281.35,    281.35,  281.35,  281.35,
  281.25,    281.25,  281.25,  281.25,
  281.1,     281.1,   281.1,   281.1,
  280.85,    280.85,  280.85,  280.85,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.6,     280.6,   280.6,   280.6,
  280.35,    280.35,  280.35,  280.35,
  279.95,    279.95,  279.95,  279.95,
  279.65,    279.65,  279.65,  279.65,
  279.4,     279.4,   279.4,   279.4,
  279.2,     279.2,   279.2,   279.2,
  279.15,    279.15,  279.15,  279.15,
  279,       279,     279,     279,
  278.9,     278.9,   278.9,   278.9,
  279.1,     279.1,   279.1,   279.1,
  279.45,    279.45,  279.45,  279.45,
  280,       280,     280,     280,
  280.75,    280.75,  280.75,  280.75,
  281.6,     281.6,   281.6,   281.6,
  282.45,    282.45,  282.45,  282.45,
  283.2,     283.2,   283.2,   283.2,
  283.85,    283.85,  283.85,  283.85,
  284.45,    284.45,  284.45,  284.45,
  284.85,    284.85,  284.85,  284.85,
  284.95,    284.95,  284.95,  284.95,
  285.25,    285.25,  285.25,  285.25,
  285.45,    285.45,  285.45,  285.45,
  285.25,    285.25,  285.25,  285.25,
  285.15,    285.15,  285.15,  285.15,
  285.2,     285.2,   285.2,   285.2,
  285.35,    285.35,  285.35,  285.35,
  285.4,     285.4,   285.4,   285.4,
  285.25,    285.25,  285.25,  285.25,
  284.9,     284.9,   284.9,   284.9,
  284.35,    284.35,  284.35,  284.35,
  283.8,     283.8,   283.8,   283.8,
  283.2,     283.2,   283.2,   283.2,
  282.55,    282.55,  282.55,  282.55,
  282.05,    282.05,  282.05,  282.05,
  281.6,     281.6,   281.6,   281.6,
  281.2,     281.2,   281.2,   281.2,
  280.95,    280.95,  280.95,  280.95,
  280.75,    280.75,  280.75,  280.75,
  280.75,    280.75,  280.75,  280.75,
  280.85,    280.85,  280.85,  280.85,
  280.6,     280.6,   280.6,   280.6,
  280.35,    280.35,  280.35,  280.35,
  280.25,    280.25,  280.25,  280.25,
  280.2,     280.2,   280.2,   280.2,
  280.2,     280.2,   280.2,   280.2,
  280.1,     280.1,   280.1,   280.1,
  280,       280,     280,     280,
  279.95,    279.95,  279.95,  279.95,
  279.9,     279.9,   279.9,   279.9,
  279.8,     279.8,   279.8,   279.8,
  279.65,    279.65,  279.65,  279.65,
  279.45,    279.45,  279.45,  279.45,
  279.35,    279.35,  279.35,  279.35,
  279.35,    279.35,  279.35,  279.35,
  279.25,    279.25,  279.25,  279.25,
  279.15,    279.15,  279.15,  279.15,
  279.15,    279.15,  279.15,  279.15,
  279.15,    279.15,  279.15,  279.15,
  279.15,    279.15,  279.15,  279.15,
  279.15,    279.15,  279.15,  279.15,
  279.2,     279.2,   279.2,   279.2,
  279.35,    279.35,  279.35,  279.35,
  279.6,     279.6,   279.6,   279.6,
  280.05,    280.05,  280.05,  280.05,
  280.8,     280.8,   280.8,   280.8,
  281.75,    281.75,  281.75,  281.75,
  282.75,    282.75,  282.75,  282.75,
  283.85,    283.85,  283.85,  283.85,
  284.8,     284.8,   284.8,   284.8,
  285.5,     285.5,   285.5,   285.5,
  285.95,    285.95,  285.95,  285.95,
  286.15,    286.15,  286.15,  286.15,
  286.3,     286.3,   286.3,   286.3,
  286.4,     286.4,   286.4,   286.4,
  286.4,     286.4,   286.4,   286.4,
  286.2,     286.2,   286.2,   286.2,
  285.85,    285.85,  285.85,  285.85,
  285.25,    285.25,  285.25,  285.25,
  284.4,     284.4,   284.4,   284.4,
  283.55,    283.55,  283.55,  283.55,
  282.85,    282.85,  282.85,  282.85,
  282.3,     282.3,   282.3,   282.3,
  281.95,    281.95,  281.95,  281.95,
  281.75,    281.75,  281.75,  281.75,
  281.55,    281.55,  281.55,  281.55,
  281.25,    281.25,  281.25,  281.25,
  280.95,    280.95,  280.95,  280.95,
  280.85,    280.85,  280.85,  280.85,
  280.75,    280.75,  280.75,  280.75,
  280.55,    280.55,  280.55,  280.55,
  280.3,     280.3,   280.3,   280.3,
  280,       280,     280,     280,
  279.75,    279.75,  279.75,  279.75,
  279.65,    279.65,  279.65,  279.65,
  279.65,    279.65,  279.65,  279.65,
  279.6,     279.6,   279.6,   279.6,
  279.55,    279.55,  279.55,  279.55,
  279.35,    279.35,  279.35,  279.35,
  278.9,     278.9,   278.9,   278.9,
  278.5,     278.5,   278.5,   278.5,
  278.2,     278.2,   278.2,   278.2,
  277.9,     277.9,   277.9,   277.9,
  277.6,     277.6,   277.6,   277.6,
  277.3,     277.3,   277.3,   277.3,
  277.25,    277.25,  277.25,  277.25,
  277.75,    277.75,  277.75,  277.75,
  278.75,    278.75,  278.75,  278.75,
  280.25,    280.25,  280.25,  280.25,
  282.05,    282.05,  282.05,  282.05,
  283.7,     283.7,   283.7,   283.7,
  285,       285,     285,     285,
  286.05,    286.05,  286.05,  286.05,
  286.95,    286.95,  286.95,  286.95,
  287.8,     287.8,   287.8,   287.8,
  288.55,    288.55,  288.55,  288.55,
  289.05,    289.05,  289.05,  289.05,
  289.2,     289.2,   289.2,   289.2,
  289.2,     289.2,   289.2,   289.2,
  289.4,     289.4,   289.4,   289.4,
  289.8,     289.8,   289.8,   289.8,
  290.35,    290.35,  290.35,  290.35,
  290.45,    290.45,  290.45,  290.45,
  290.15,    290.15,  290.15,  290.15,
  289.9,     289.9,   289.9,   289.9,
  289.3,     289.3,   289.3,   289.3,
  288.35,    288.35,  288.35,  288.35,
  287.1,     287.1,   287.1,   287.1,
  285.65,    285.65,  285.65,  285.65,
  284.4,     284.4,   284.4,   284.4,
  283.5,     283.5,   283.5,   283.5,
  282.75,    282.75,  282.75,  282.75,
  281.9,     281.9,   281.9,   281.9,
  280.85,    280.85,  280.85,  280.85,
  279.75,    279.75,  279.75,  279.75,
  278.9,     278.9,   278.9,   278.9,
  278.4,     278.4,   278.4,   278.4,
  278.1,     278.1,   278.1,   278.1,
  277.9,     277.9,   277.9,   277.9,
  277.65,    277.65,  277.65,  277.65,
  277.35,    277.35,  277.35,  277.35,
  277.15,    277.15,  277.15,  277.15,
  276.9,     276.9,   276.9,   276.9,
  276.75,    276.75,  276.75,  276.75,
  276.75,    276.75,  276.75,  276.75,
  276.75,    276.75,  276.75,  276.75,
  276.7,     276.7,   276.7,   276.7,
  276.7,     276.7,   276.7,   276.7,
  276.8,     276.8,   276.8,   276.8,
  276.85,    276.85,  276.85,  276.85,
  276.75,    276.75,  276.75,  276.75,
  276.5,     276.5,   276.5,   276.5,
  276.4,     276.4,   276.4,   276.4,
  276.45,    276.45,  276.45,  276.45,
  276.45,    276.45,  276.45,  276.45,
  276.45,    276.45,  276.45,  276.45,
  276.5,     276.5,   276.5,   276.5,
  276.75,    276.75,  276.75,  276.75,
  277.1,     277.1,   277.1,   277.1,
  277.45,    277.45,  277.45,  277.45,
  277.8,     277.8,   277.8,   277.8,
  278.2,     278.2,   278.2,   278.2,
  278.65,    278.65,  278.65,  278.65,
  279.1,     279.1,   279.1,   279.1,
  279.85,    279.85,  279.85,  279.85,
  280.75,    280.75,  280.75,  280.75,
  281.45,    281.45,  281.45,  281.45,
  282.1,     282.1,   282.1,   282.1,
  282.55,    282.55,  282.55,  282.55,
  282.25,    282.25,  282.25,  282.25,
  281.4,     281.4,   281.4,   281.4,
  280.7,     280.7,   280.7,   280.7,
  280.25,    280.25,  280.25,  280.25,
  279.8,     279.8,   279.8,   279.8,
  279.4,     279.4,   279.4,   279.4,
  279.05,    279.05,  279.05,  279.05,
  278.6,     278.6,   278.6,   278.6,
  278.1,     278.1,   278.1,   278.1,
  277.8,     277.8,   277.8,   277.8,
  277.55,    277.55,  277.55,  277.55,
  277.3,     277.3,   277.3,   277.3,
  277.25,    277.25,  277.25,  277.25,
  277.25,    277.25,  277.25,  277.25,
  277.25,    277.25,  277.25,  277.25,
  277.25,    277.25,  277.25,  277.25,
  277.25,    277.25,  277.25,  277.25,
  277.2,     277.2,   277.2,   277.2,
  277.1,     277.1,   277.1,   277.1,
  276.95,    276.95,  276.95,  276.95,
  276.8,     276.8,   276.8,   276.8,
  276.65,    276.65,  276.65,  276.65,
  276.5,     276.5,   276.5,   276.5,
  276.4,     276.4,   276.4,   276.4,
  276.3,     276.3,   276.3,   276.3,
  276.15,    276.15,  276.15,  276.15,
  276.05,    276.05,  276.05,  276.05,
  276,       276,     276,     276,
  275.85,    275.85,  275.85,  275.85,
  275.75,    275.75,  275.75,  275.75,
  275.7,     275.7,   275.7,   275.7,
  275.6,     275.6,   275.6,   275.6,
  275.55,    275.55,  275.55,  275.55,
  275.6,     275.6,   275.6,   275.6,
  275.7,     275.7,   275.7,   275.7,
  275.8,     275.8,   275.8,   275.8,
  276.1,     276.1,   276.1,   276.1,
  276.55,    276.55,  276.55,  276.55,
  277.05,    277.05,  277.05,  277.05,
  278,       278,     278,     278,
  279.45,    279.45,  279.45,  279.45,
  281.05,    281.05,  281.05,  281.05,
  282.25,    282.25,  282.25,  282.25,
  283.1,     283.1,   283.1,   283.1,
  283.65,    283.65,  283.65,  283.65,
  284.15,    284.15,  284.15,  284.15,
  284.9,     284.9,   284.9,   284.9,
  285.55,    285.55,  285.55,  285.55,
  286.1,     286.1,   286.1,   286.1,
  286.2,     286.2,   286.2,   286.2,
  285.9,     285.9,   285.9,   285.9,
  285.7,     285.7,   285.7,   285.7,
  285.4,     285.4,   285.4,   285.4,
  284.8,     284.8,   284.8,   284.8,
  284.25,    284.25,  284.25,  284.25,
  283.8,     283.8,   283.8,   283.8,
  283.4,     283.4,   283.4,   283.4,
  282.95,    282.95,  282.95,  282.95,
  282.45,    282.45,  282.45,  282.45,
  281.95,    281.95,  281.95,  281.95,
  281.55,    281.55,  281.55,  281.55,
  281.2,     281.2,   281.2,   281.2,
  280.8,     280.8,   280.8,   280.8,
  280.5,     280.5,   280.5,   280.5,
  280.15,    280.15,  280.15,  280.15,
  280.05,    280.05,  280.05,  280.05,
  280.25,    280.25,  280.25,  280.25,
  280.15,    280.15,  280.15,  280.15,
  279.75,    279.75,  279.75,  279.75,
  279.5,     279.5,   279.5,   279.5,
  279.5,     279.5,   279.5,   279.5,
  279.75,    279.75,  279.75,  279.75,
  280.15,    280.15,  280.15,  280.15,
  280.5,     280.5,   280.5,   280.5,
  280.7,     280.7,   280.7,   280.7,
  280.8,     280.8,   280.8,   280.8,
  280.9,     280.9,   280.9,   280.9,
  280.8,     280.8,   280.8,   280.8,
  280.4,     280.4,   280.4,   280.4,
  280.05,    280.05,  280.05,  280.05,
  279.95,    279.95,  279.95,  279.95,
  280.1,     280.1,   280.1,   280.1,
  280.65,    280.65,  280.65,  280.65,
  281.5,     281.5,   281.5,   281.5,
  282.25,    282.25,  282.25,  282.25,
  283.05,    283.05,  283.05,  283.05,
  283.9,     283.9,   283.9,   283.9,
  284.5,     284.5,   284.5,   284.5,
  285.1,     285.1,   285.1,   285.1,
  285.75,    285.75,  285.75,  285.75,
  286.35,    286.35,  286.35,  286.35,
  286.7,     286.7,   286.7,   286.7,
  286.65,    286.65,  286.65,  286.65,
  286.75,    286.75,  286.75,  286.75,
  287.2,     287.2,   287.2,   287.2,
  287.15,    287.15,  287.15,  287.15,
  286.8,     286.8,   286.8,   286.8,
  286.65,    286.65,  286.65,  286.65,
  286.5,     286.5,   286.5,   286.5,
  286.25,    286.25,  286.25,  286.25,
  285.65,    285.65,  285.65,  285.65,
  284.3,     284.3,   284.3,   284.3,
  283.1,     283.1,   283.1,   283.1,
  282.8,     282.8,   282.8,   282.8,
  282.5,     282.5,   282.5,   282.5,
  282,       282,     282,     282,
  281.65,    281.65,  281.65,  281.65,
  281.55,    281.55,  281.55,  281.55,
  281.55,    281.55,  281.55,  281.55,
  281.5,     281.5,   281.5,   281.5,
  281.45,    281.45,  281.45,  281.45,
  281.45,    281.45,  281.45,  281.45,
  281.45,    281.45,  281.45,  281.45,
  281.4,     281.4,   281.4,   281.4,
  281.25,    281.25,  281.25,  281.25,
  281.05,    281.05,  281.05,  281.05,
  280.8,     280.8,   280.8,   280.8,
  280.65,    280.65,  280.65,  280.65,
  280.6,     280.6,   280.6,   280.6,
  280.55,    280.55,  280.55,  280.55,
  280.5,     280.5,   280.5,   280.5,
  280.4,     280.4,   280.4,   280.4,
  280.4,     280.4,   280.4,   280.4,
  280.45,    280.45,  280.45,  280.45,
  280.45,    280.45,  280.45,  280.45,
  280.45,    280.45,  280.45,  280.45,
  280.5,     280.5,   280.5,   280.5,
  280.6,     280.6,   280.6,   280.6,
  280.7,     280.7,   280.7,   280.7,
  280.8,     280.8,   280.8,   280.8,
  280.95,    280.95,  280.95,  280.95,
  281.15,    281.15,  281.15,  281.15,
  281.35,    281.35,  281.35,  281.35,
  281.5,     281.5,   281.5,   281.5,
  281.55,    281.55,  281.55,  281.55,
  281.45,    281.45,  281.45,  281.45,
  281.3,     281.3,   281.3,   281.3,
  281.3,     281.3,   281.3,   281.3,
  281.45,    281.45,  281.45,  281.45,
  281.65,    281.65,  281.65,  281.65,
  281.85,    281.85,  281.85,  281.85,
  282,       282,     282,     282,
  282.05,    282.05,  282.05,  282.05,
  282.15,    282.15,  282.15,  282.15,
  282.2,     282.2,   282.2,   282.2,
  282.15,    282.15,  282.15,  282.15,
  282.15,    282.15,  282.15,  282.15,
  282.2,     282.2,   282.2,   282.2,
  282.3,     282.3,   282.3,   282.3,
  282.35,    282.35,  282.35,  282.35,
  282.35,    282.35,  282.35,  282.35,
  282.35,    282.35,  282.35,  282.35,
  282.35,    282.35,  282.35,  282.35,
  282.25,    282.25,  282.25,  282.25,
  281.95,    281.95,  281.95,  281.95,
  281.7,     281.7,   281.7,   281.7,
  281.65,    281.65,  281.65,  281.65,
  281.6,     281.6,   281.6,   281.6,
  281.55,    281.55,  281.55,  281.55,
  281.6,     281.6,   281.6,   281.6,
  281.55,    281.55,  281.55,  281.55,
  281.3,     281.3,   281.3,   281.3,
  281.1,     281.1,   281.1,   281.1,
  281.15,    281.15,  281.15,  281.15,
  281.35,    281.35,  281.35,  281.35,
  281.35,    281.35,  281.35,  281.35,
  281.3,     281.3,   281.3,   281.3,
  281.45,    281.45,  281.45,  281.45,
  281.5,     281.5,   281.5,   281.5,
  281.4,     281.4,   281.4,   281.4,
  281.35,    281.35,  281.35,  281.35,
  281.4,     281.4,   281.4,   281.4,
  281.5,     281.5,   281.5,   281.5,
  281.55,    281.55,  281.55,  281.55,
  281.5,     281.5,   281.5,   281.5,
  281.5,     281.5,   281.5,   281.5,
  281.6,     281.6,   281.6,   281.6,
  281.7,     281.7,   281.7,   281.7,
  281.9,     281.9,   281.9,   281.9,
  282.25,    282.25,  282.25,  282.25,
  282.55,    282.55,  282.55,  282.55,
  282.7,     282.7,   282.7,   282.7,
  282.9,     282.9,   282.9,   282.9,
  283.15,    283.15,  283.15,  283.15,
  283.25,    283.25,  283.25,  283.25,
  282.95,    282.95,  282.95,  282.95,
  282.3,     282.3,   282.3,   282.3,
  281.9,     281.9,   281.9,   281.9,
  281.85,    281.85,  281.85,  281.85,
  281.95,    281.95,  281.95,  281.95,
  282.15,    282.15,  282.15,  282.15,
  282.35,    282.35,  282.35,  282.35,
  282.5,     282.5,   282.5,   282.5,
  282.6,     282.6,   282.6,   282.6,
  282.7,     282.7,   282.7,   282.7,
  282.7,     282.7,   282.7,   282.7,
  282.6,     282.6,   282.6,   282.6,
  282.55,    282.55,  282.55,  282.55,
  282.5,     282.5,   282.5,   282.5,
  282.45,    282.45,  282.45,  282.45,
  282.5,     282.5,   282.5,   282.5,
  282.5,     282.5,   282.5,   282.5,
  282.45,    282.45,  282.45,  282.45,
  282.4,     282.4,   282.4,   282.4,
  282.35,    282.35,  282.35,  282.35,
  282.35,    282.35,  282.35,  282.35,
  282.35,    282.35,  282.35,  282.35,
  282.3,     282.3,   282.3,   282.3,
  282,       282,     282,     282,
  281.65,    281.65,  281.65,  281.65,
  281.45,    281.45,  281.45,  281.45,
  281.3,     281.3,   281.3,   281.3,
  281.2,     281.2,   281.2,   281.2,
  281,       281,     281,     281,
  280.75,    280.75,  280.75,  280.75,
  280.6,     280.6,   280.6,   280.6,
  280.55,    280.55,  280.55,  280.55,
  280.55,    280.55,  280.55,  280.55,
  280.5,     280.5,   280.5,   280.5,
  280.5,     280.5,   280.5,   280.5,
  280.55,    280.55,  280.55,  280.55,
  280.55,    280.55,  280.55,  280.55,
  280.6,     280.6,   280.6,   280.6,
  280.75,    280.75,  280.75,  280.75,
  280.95,    280.95,  280.95,  280.95,
  281.1,     281.1,   281.1,   281.1,
  281.2,     281.2,   281.2,   281.2,
  281.35,    281.35,  281.35,  281.35,
  281.55,    281.55,  281.55,  281.55,
  281.9,     281.9,   281.9,   281.9,
  282.4,     282.4,   282.4,   282.4,
  282.8,     282.8,   282.8,   282.8,
  283,       283,     283,     283,
  283.1,     283.1,   283.1,   283.1,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  283.1,     283.1,   283.1,   283.1,
  283,       283,     283,     283,
  282.9,     282.9,   282.9,   282.9,
  282.95,    282.95,  282.95,  282.95,
  283.05,    283.05,  283.05,  283.05,
  283.1,     283.1,   283.1,   283.1,
  283.15,    283.15,  283.15,  283.15,
  282.9,     282.9,   282.9,   282.9,
  282.5,     282.5,   282.5,   282.5,
  282.3,     282.3,   282.3,   282.3,
  282.25,    282.25,  282.25,  282.25,
  282.25,    282.25,  282.25,  282.25,
  282.2,     282.2,   282.2,   282.2,
  282.2,     282.2,   282.2,   282.2,
  282.25,    282.25,  282.25,  282.25,
  282.25,    282.25,  282.25,  282.25,
  282.25,    282.25,  282.25,  282.25,
  282.3,     282.3,   282.3,   282.3,
  282.25,    282.25,  282.25,  282.25,
  281.8,     281.8,   281.8,   281.8,
  281.45,    281.45,  281.45,  281.45,
  281.6,     281.6,   281.6,   281.6,
  281.85,    281.85,  281.85,  281.85,
  282.05,    282.05,  282.05,  282.05,
  282.4,     282.4,   282.4,   282.4,
  282.6,     282.6,   282.6,   282.6,
  282.55,    282.55,  282.55,  282.55,
  282.45,    282.45,  282.45,  282.45,
  282.25,    282.25,  282.25,  282.25,
  282.1,     282.1,   282.1,   282.1,
  281.95,    281.95,  281.95,  281.95,
  281.75,    281.75,  281.75,  281.75,
  281.55,    281.55,  281.55,  281.55,
  281.35,    281.35,  281.35,  281.35,
  281.15,    281.15,  281.15,  281.15,
  280.9,     280.9,   280.9,   280.9,
  280.7,     280.7,   280.7,   280.7,
  280.7,     280.7,   280.7,   280.7,
  281,       281,     281,     281,
  281.3,     281.3,   281.3,   281.3,
  281.5,     281.5,   281.5,   281.5,
  281.7,     281.7,   281.7,   281.7,
  281.75,    281.75,  281.75,  281.75,
  281.85,    281.85,  281.85,  281.85,
  282.2,     282.2,   282.2,   282.2,
  282.5,     282.5,   282.5,   282.5,
  282.65,    282.65,  282.65,  282.65,
  283,       283,     283,     283,
  283.4,     283.4,   283.4,   283.4,
  283.45,    283.45,  283.45,  283.45,
  283.45,    283.45,  283.45,  283.45,
  283.65,    283.65,  283.65,  283.65,
  283.55,    283.55,  283.55,  283.55,
  283.05,    283.05,  283.05,  283.05,
  282.65,    282.65,  282.65,  282.65,
  282.3,     282.3,   282.3,   282.3,
  281.9,     281.9,   281.9,   281.9,
  281.6,     281.6,   281.6,   281.6,
  281.1,     281.1,   281.1,   281.1,
  280.45,    280.45,  280.45,  280.45,
  280.05,    280.05,  280.05,  280.05,
  279.75,    279.75,  279.75,  279.75,
  279.4,     279.4,   279.4,   279.4,
  279.15,    279.15,  279.15,  279.15,
  278.9,     278.9,   278.9,   278.9,
  278.5,     278.5,   278.5,   278.5,
  278.05,    278.05,  278.05,  278.05,
  277.7,     277.7,   277.7,   277.7,
  277.4,     277.4,   277.4,   277.4,
  277.15,    277.15,  277.15,  277.15,
  276.95,    276.95,  276.95,  276.95,
  276.85,    276.85,  276.85,  276.85,
  276.75,    276.75,  276.75,  276.75,
  276.6,     276.6,   276.6,   276.6,
  276.7,     276.7,   276.7,   276.7,
  277,       277,     277,     277,
  277.15,    277.15,  277.15,  277.15,
  277.3,     277.3,   277.3,   277.3,
  277.5,     277.5,   277.5,   277.5,
  277.6,     277.6,   277.6,   277.6,
  277.75,    277.75,  277.75,  277.75,
  277.95,    277.95,  277.95,  277.95,
  278.1,     278.1,   278.1,   278.1,
  278.3,     278.3,   278.3,   278.3,
  278.6,     278.6,   278.6,   278.6,
  278.9,     278.9,   278.9,   278.9,
  279.25,    279.25,  279.25,  279.25,
  279.6,     279.6,   279.6,   279.6,
  279.85,    279.85,  279.85,  279.85,
  280.35,    280.35,  280.35,  280.35,
  281.15,    281.15,  281.15,  281.15,
  281.7,     281.7,   281.7,   281.7,
  282.1,     282.1,   282.1,   282.1,
  282.6,     282.6,   282.6,   282.6,
  282.9,     282.9,   282.9,   282.9,
  282.2,     282.2,   282.2,   282.2,
  281.25,    281.25,  281.25,  281.25,
  281.05,    281.05,  281.05,  281.05,
  281.1,     281.1,   281.1,   281.1,
  281.3,     281.3,   281.3,   281.3,
  281.25,    281.25,  281.25,  281.25,
  280.7,     280.7,   280.7,   280.7,
  280.25,    280.25,  280.25,  280.25,
  280.15,    280.15,  280.15,  280.15,
  280.2,     280.2,   280.2,   280.2,
  280.25,    280.25,  280.25,  280.25,
  280.25,    280.25,  280.25,  280.25,
  279.15,    279.15,  279.15,  279.15,
  278,       278,     278,     278,
  277.8,     277.8,   277.8,   277.8,
  277.65,    277.65,  277.65,  277.65,
  277.6,     277.6,   277.6,   277.6,
  277.6,     277.6,   277.6,   277.6,
  277.75,    277.75,  277.75,  277.75,
  278.1,     278.1,   278.1,   278.1,
  278.55,    278.55,  278.55,  278.55,
  278.6,     278.6,   278.6,   278.6,
  278.65,    278.65,  278.65,  278.65,
  278.95,    278.95,  278.95,  278.95,
  279.3,     279.3,   279.3,   279.3,
  279.65,    279.65,  279.65,  279.65,
  279.75,    279.75,  279.75,  279.75,
  279.55,    279.55,  279.55,  279.55,
  279.3,     279.3,   279.3,   279.3,
  279.3,     279.3,   279.3,   279.3,
  279.5,     279.5,   279.5,   279.5,
  279.45,    279.45,  279.45,  279.45,
  279.15,    279.15,  279.15,  279.15,
  279,       279,     279,     279,
  278.95,    278.95,  278.95,  278.95,
  279.05,    279.05,  279.05,  279.05,
  279.2,     279.2,   279.2,   279.2,
  279.3,     279.3,   279.3,   279.3,
  279.35,    279.35,  279.35,  279.35,
  279.45,    279.45,  279.45,  279.45,
  279.6,     279.6,   279.6,   279.6,
  279.65,    279.65,  279.65,  279.65,
  279.6,     279.6,   279.6,   279.6,
  279.65,    279.65,  279.65,  279.65,
  280,       280,     280,     280,
  280.45,    280.45,  280.45,  280.45,
  280.7,     280.7,   280.7,   280.7,
  280.7,     280.7,   280.7,   280.7,
  280.7,     280.7,   280.7,   280.7,
  281,       281,     281,     281,
  281.2,     281.2,   281.2,   281.2,
  280.8,     280.8,   280.8,   280.8,
  280.3,     280.3,   280.3,   280.3,
  280.05,    280.05,  280.05,  280.05,
  279.7,     279.7,   279.7,   279.7,
  279.05,    279.05,  279.05,  279.05,
  278.25,    278.25,  278.25,  278.25,
  277.6,     277.6,   277.6,   277.6,
  277.2,     277.2,   277.2,   277.2,
  277,       277,     277,     277,
  276.85,    276.85,  276.85,  276.85,
  276.7,     276.7,   276.7,   276.7,
  276.55,    276.55,  276.55,  276.55,
  276.4,     276.4,   276.4,   276.4,
  276.25,    276.25,  276.25,  276.25,
  276.1,     276.1,   276.1,   276.1,
  276.05,    276.05,  276.05,  276.05,
  276,       276,     276,     276,
  275.9,     275.9,   275.9,   275.9,
  275.8,     275.8,   275.8,   275.8,
  275.75,    275.75,  275.75,  275.75,
  275.7,     275.7,   275.7,   275.7,
  275.6,     275.6,   275.6,   275.6,
  275.5,     275.5,   275.5,   275.5,
  275.4,     275.4,   275.4,   275.4,
  275.25,    275.25,  275.25,  275.25,
  275.15,    275.15,  275.15,  275.15,
  275.05,    275.05,  275.05,  275.05,
  274.9,     274.9,   274.9,   274.9,
  274.8,     274.8,   274.8,   274.8,
  274.7,     274.7,   274.7,   274.7,
  274.5,     274.5,   274.5,   274.5,
  274.4,     274.4,   274.4,   274.4,
  274.45,    274.45,  274.45,  274.45,
  274.4,     274.4,   274.4,   274.4,
  274.55,    274.55,  274.55,  274.55,
  275.05,    275.05,  275.05,  275.05,
  275.6,     275.6,   275.6,   275.6,
  275.9,     275.9,   275.9,   275.9,
  276.1,     276.1,   276.1,   276.1,
  276.45,    276.45,  276.45,  276.45,
  276.8,     276.8,   276.8,   276.8,
  277.2,     277.2,   277.2,   277.2,
  277.7,     277.7,   277.7,   277.7,
  278.25,    278.25,  278.25,  278.25,
  278.55,    278.55,  278.55,  278.55,
  278.45,    278.45,  278.45,  278.45,
  278.3,     278.3,   278.3,   278.3,
  278.2,     278.2,   278.2,   278.2,
  278.4,     278.4,   278.4,   278.4,
  278.7,     278.7,   278.7,   278.7,
  278.85,    278.85,  278.85,  278.85,
  278.95,    278.95,  278.95,  278.95,
  278.8,     278.8,   278.8,   278.8,
  278.45,    278.45,  278.45,  278.45,
  278.15,    278.15,  278.15,  278.15,
  278.15,    278.15,  278.15,  278.15,
  278.3,     278.3,   278.3,   278.3,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.3,     278.3,   278.3,   278.3,
  278.25,    278.25,  278.25,  278.25,
  278.25,    278.25,  278.25,  278.25,
  278.2,     278.2,   278.2,   278.2,
  278.2,     278.2,   278.2,   278.2,
  278.3,     278.3,   278.3,   278.3,
  278.15,    278.15,  278.15,  278.15,
  277.65,    277.65,  277.65,  277.65,
  277.15,    277.15,  277.15,  277.15,
  277,       277,     277,     277,
  277.15,    277.15,  277.15,  277.15,
  277.3,     277.3,   277.3,   277.3,
  277.45,    277.45,  277.45,  277.45,
  277.55,    277.55,  277.55,  277.55,
  277.55,    277.55,  277.55,  277.55,
  277.45,    277.45,  277.45,  277.45,
  277.35,    277.35,  277.35,  277.35,
  277.45,    277.45,  277.45,  277.45,
  277.55,    277.55,  277.55,  277.55,
  277.6,     277.6,   277.6,   277.6,
  277.35,    277.35,  277.35,  277.35,
  276.85,    276.85,  276.85,  276.85,
  276.8,     276.8,   276.8,   276.8,
  277.15,    277.15,  277.15,  277.15,
  277.6,     277.6,   277.6,   277.6,
  278.05,    278.05,  278.05,  278.05,
  278.45,    278.45,  278.45,  278.45,
  278.9,     278.9,   278.9,   278.9,
  279.25,    279.25,  279.25,  279.25,
  279.2,     279.2,   279.2,   279.2,
  279.15,    279.15,  279.15,  279.15,
  279.3,     279.3,   279.3,   279.3,
  279.45,    279.45,  279.45,  279.45,
  279.6,     279.6,   279.6,   279.6,
  279.9,     279.9,   279.9,   279.9,
  280.05,    280.05,  280.05,  280.05,
  279.7,     279.7,   279.7,   279.7,
  279.85,    279.85,  279.85,  279.85,
  280.45,    280.45,  280.45,  280.45,
  280.75,    280.75,  280.75,  280.75,
  280.5,     280.5,   280.5,   280.5,
  280.05,    280.05,  280.05,  280.05,
  279.85,    279.85,  279.85,  279.85,
  279.25,    279.25,  279.25,  279.25,
  278.55,    278.55,  278.55,  278.55,
  278.2,     278.2,   278.2,   278.2,
  277.85,    277.85,  277.85,  277.85,
  277.25,    277.25,  277.25,  277.25,
  276.5,     276.5,   276.5,   276.5,
  276,       276,     276,     276,
  275.45,    275.45,  275.45,  275.45,
  274.75,    274.75,  274.75,  274.75,
  274.4,     274.4,   274.4,   274.4,
  274.25,    274.25,  274.25,  274.25,
  274.1,     274.1,   274.1,   274.1,
  273.9,     273.9,   273.9,   273.9,
  273.6,     273.6,   273.6,   273.6,
  273.4,     273.4,   273.4,   273.4,
  272.95,    272.95,  272.95,  272.95,
  272.7,     272.7,   272.7,   272.7,
  272.85,    272.85,  272.85,  272.85,
  272.7,     272.7,   272.7,   272.7,
  272.5,     272.5,   272.5,   272.5,
  272.3,     272.3,   272.3,   272.3,
  272.1,     272.1,   272.1,   272.1,
  271.85,    271.85,  271.85,  271.85,
  271.4,     271.4,   271.4,   271.4,
  271.4,     271.4,   271.4,   271.4,
  271.75,    271.75,  271.75,  271.75,
  271.25,    271.25,  271.25,  271.25,
  270.65,    270.65,  270.65,  270.65,
  270.95,    270.95,  270.95,  270.95,
  271.6,     271.6,   271.6,   271.6,
  272.4,     272.4,   272.4,   272.4,
  273.6,     273.6,   273.6,   273.6,
  275.5,     275.5,   275.5,   275.5,
  277.1,     277.1,   277.1,   277.1,
  277.6,     277.6,   277.6,   277.6,
  277.9,     277.9,   277.9,   277.9,
  278.4,     278.4,   278.4,   278.4,
  278.8,     278.8,   278.8,   278.8,
  279.1,     279.1,   279.1,   279.1,
  279.25,    279.25,  279.25,  279.25,
  279.65,    279.65,  279.65,  279.65,
  279.95,    279.95,  279.95,  279.95,
  280.15,    280.15,  280.15,  280.15,
  280.5,     280.5,   280.5,   280.5,
  280.65,    280.65,  280.65,  280.65,
  280.75,    280.75,  280.75,  280.75,
  280.85,    280.85,  280.85,  280.85,
  280.85,    280.85,  280.85,  280.85,
  280.6,     280.6,   280.6,   280.6,
  280.2,     280.2,   280.2,   280.2,
  279.6,     279.6,   279.6,   279.6,
  279.1,     279.1,   279.1,   279.1,
  278.65,    278.65,  278.65,  278.65,
  278.3,     278.3,   278.3,   278.3,
  278.2,     278.2,   278.2,   278.2,
  278.1,     278.1,   278.1,   278.1,
  278,       278,     278,     278,
  277.9,     277.9,   277.9,   277.9,
  277.85,    277.85,  277.85,  277.85,
  277.9,     277.9,   277.9,   277.9,
  278,       278,     278,     278,
  278,       278,     278,     278,
  277.95,    277.95,  277.95,  277.95,
  278.05,    278.05,  278.05,  278.05,
  278.1,     278.1,   278.1,   278.1,
  277.95,    277.95,  277.95,  277.95,
  277.7,     277.7,   277.7,   277.7,
  277.5,     277.5,   277.5,   277.5,
  277.5,     277.5,   277.5,   277.5,
  277.5,     277.5,   277.5,   277.5,
  277.4,     277.4,   277.4,   277.4,
  277.45,    277.45,  277.45,  277.45,
  277.75,    277.75,  277.75,  277.75,
  278,       278,     278,     278,
  278.05,    278.05,  278.05,  278.05,
  278,       278,     278,     278,
  277.6,     277.6,   277.6,   277.6,
  277.35,    277.35,  277.35,  277.35,
  277.5,     277.5,   277.5,   277.5,
  277.65,    277.65,  277.65,  277.65,
  277.9,     277.9,   277.9,   277.9,
  277.95,    277.95,  277.95,  277.95,
  277.75,    277.75,  277.75,  277.75,
  277.65,    277.65,  277.65,  277.65,
  277.6,     277.6,   277.6,   277.6,
  277.5,     277.5,   277.5,   277.5,
  277.5,     277.5,   277.5,   277.5,
  277.65,    277.65,  277.65,  277.65,
  277.8,     277.8,   277.8,   277.8,
  277.95,    277.95,  277.95,  277.95,
  278.2,     278.2,   278.2,   278.2,
  278.35,    278.35,  278.35,  278.35,
  278.4,     278.4,   278.4,   278.4,
  278.5,     278.5,   278.5,   278.5,
  278.6,     278.6,   278.6,   278.6,
  278.7,     278.7,   278.7,   278.7,
  278.8,     278.8,   278.8,   278.8,
  278.9,     278.9,   278.9,   278.9,
  278.95,    278.95,  278.95,  278.95,
  278.9,     278.9,   278.9,   278.9,
  278.8,     278.8,   278.8,   278.8,
  278.7,     278.7,   278.7,   278.7,
  278.75,    278.75,  278.75,  278.75,
  278.8,     278.8,   278.8,   278.8,
  278.8,     278.8,   278.8,   278.8,
  278.7,     278.7,   278.7,   278.7,
  278.45,    278.45,  278.45,  278.45,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.4,     278.4,   278.4,   278.4,
  278.4,     278.4,   278.4,   278.4,
  278.25,    278.25,  278.25,  278.25,
  278.1,     278.1,   278.1,   278.1,
  278,       278,     278,     278,
  277.95,    277.95,  277.95,  277.95,
  277.95,    277.95,  277.95,  277.95,
  277.95,    277.95,  277.95,  277.95,
  277.9,     277.9,   277.9,   277.9,
  277.8,     277.8,   277.8,   277.8,
  277.75,    277.75,  277.75,  277.75,
  277.65,    277.65,  277.65,  277.65,
  277.5,     277.5,   277.5,   277.5,
  277.45,    277.45,  277.45,  277.45,
  277.5,     277.5,   277.5,   277.5,
  277.6,     277.6,   277.6,   277.6,
  277.75,    277.75,  277.75,  277.75,
  277.9,     277.9,   277.9,   277.9,
  277.95,    277.95,  277.95,  277.95,
  278.05,    278.05,  278.05,  278.05,
  278.25,    278.25,  278.25,  278.25,
  278.5,     278.5,   278.5,   278.5,
  278.8,     278.8,   278.8,   278.8,
  279.1,     279.1,   279.1,   279.1,
  279.35,    279.35,  279.35,  279.35,
  279.6,     279.6,   279.6,   279.6,
  279.8,     279.8,   279.8,   279.8,
  280,       280,     280,     280,
  280.25,    280.25,  280.25,  280.25,
  280.45,    280.45,  280.45,  280.45,
  280.55,    280.55,  280.55,  280.55,
  280.55,    280.55,  280.55,  280.55,
  280.55,    280.55,  280.55,  280.55,
  280.6,     280.6,   280.6,   280.6,
  280.6,     280.6,   280.6,   280.6,
  280.45,    280.45,  280.45,  280.45,
  280.25,    280.25,  280.25,  280.25,
  280.1,     280.1,   280.1,   280.1,
  280.05,    280.05,  280.05,  280.05,
  280,       280,     280,     280,
  279.85,    279.85,  279.85,  279.85,
  279.75,    279.75,  279.75,  279.75,
  279.55,    279.55,  279.55,  279.55,
  279.35,    279.35,  279.35,  279.35,
  279.3,     279.3,   279.3,   279.3,
  279.15,    279.15,  279.15,  279.15,
  279,       279,     279,     279,
  278.95,    278.95,  278.95,  278.95,
  279,       279,     279,     279,
  279.05,    279.05,  279.05,  279.05,
  279,       279,     279,     279,
  278.95,    278.95,  278.95,  278.95,
  278.9,     278.9,   278.9,   278.9,
  278.85,    278.85,  278.85,  278.85,
  278.7,     278.7,   278.7,   278.7,
  278.5,     278.5,   278.5,   278.5,
  278.45,    278.45,  278.45,  278.45,
  278.45,    278.45,  278.45,  278.45,
  278.45,    278.45,  278.45,  278.45,
  278.4,     278.4,   278.4,   278.4,
  278.35,    278.35,  278.35,  278.35,
  278.3,     278.3,   278.3,   278.3,
  278.25,    278.25,  278.25,  278.25,
  278.3,     278.3,   278.3,   278.3,
  278.4,     278.4,   278.4,   278.4,
  278.55,    278.55,  278.55,  278.55,
  278.75,    278.75,  278.75,  278.75,
  279.05,    279.05,  279.05,  279.05,
  279.5,     279.5,   279.5,   279.5,
  279.85,    279.85,  279.85,  279.85,
  280.15,    280.15,  280.15,  280.15,
  280.45,    280.45,  280.45,  280.45,
  280.75,    280.75,  280.75,  280.75,
  280.9,     280.9,   280.9,   280.9,
  280.9,     280.9,   280.9,   280.9,
  281.1,     281.1,   281.1,   281.1,
  281.4,     281.4,   281.4,   281.4,
  281.65,    281.65,  281.65,  281.65,
  281.85,    281.85,  281.85,  281.85,
  282.1,     282.1,   282.1,   282.1,
  282.25,    282.25,  282.25,  282.25,
  282.25,    282.25,  282.25,  282.25,
  282.15,    282.15,  282.15,  282.15,
  282.1,     282.1,   282.1,   282.1,
  282.1,     282.1,   282.1,   282.1,
  281.95,    281.95,  281.95,  281.95,
  281.75,    281.75,  281.75,  281.75,
  281.4,     281.4,   281.4,   281.4,
  281.1,     281.1,   281.1,   281.1,
  281,       281,     281,     281,
  280.5,     280.5,   280.5,   280.5,
  279.75,    279.75,  279.75,  279.75,
  279.35,    279.35,  279.35,  279.35,
  279.2,     279.2,   279.2,   279.2,
  279,       279,     279,     279,
  278.7,     278.7,   278.7,   278.7,
  278.45,    278.45,  278.45,  278.45,
  278.15,    278.15,  278.15,  278.15,
  277.8,     277.8,   277.8,   277.8,
  277.65,    277.65,  277.65,  277.65,
  277.4,     277.4,   277.4,   277.4,
  276.9,     276.9,   276.9,   276.9,
  276.75,    276.75,  276.75,  276.75,
  276.85,    276.85,  276.85,  276.85,
  277.1,     277.1,   277.1,   277.1,
  277.65,    277.65,  277.65,  277.65,
  278.15,    278.15,  278.15,  278.15,
  278.35,    278.35,  278.35,  278.35,
  278.45,    278.45,  278.45,  278.45,
  278.65,    278.65,  278.65,  278.65,
  278.95,    278.95,  278.95,  278.95,
  279.55,    279.55,  279.55,  279.55,
  280.25,    280.25,  280.25,  280.25,
  280.75,    280.75,  280.75,  280.75,
  281.1,     281.1,   281.1,   281.1,
  281.4,     281.4,   281.4,   281.4,
  281.75,    281.75,  281.75,  281.75,
  282.25,    282.25,  282.25,  282.25,
  282.55,    282.55,  282.55,  282.55,
  282.6,     282.6,   282.6,   282.6,
  282.8,     282.8,   282.8,   282.8,
  283.35,    283.35,  283.35,  283.35,
  283.9,     283.9,   283.9,   283.9,
  284.3,     284.3,   284.3,   284.3,
  284.65,    284.65,  284.65,  284.65,
  284.85,    284.85,  284.85,  284.85,
  285.05,    285.05,  285.05,  285.05,
  285.2,     285.2,   285.2,   285.2,
  285.35,    285.35,  285.35,  285.35,
  285.45,    285.45,  285.45,  285.45,
  285.5,     285.5,   285.5,   285.5,
  285.55,    285.55,  285.55,  285.55,
  285.6,     285.6,   285.6,   285.6,
  285.6,     285.6,   285.6,   285.6,
  285.4,     285.4,   285.4,   285.4,
  284.65,    284.65,  284.65,  284.65,
  283.55,    283.55,  283.55,  283.55,
  283,       283,     283,     283,
  282.95,    282.95,  282.95,  282.95,
  283.05,    283.05,  283.05,  283.05,
  283.25,    283.25,  283.25,  283.25,
  283.4,     283.4,   283.4,   283.4,
  283.5,     283.5,   283.5,   283.5,
  283.6,     283.6,   283.6,   283.6,
  283.75,    283.75,  283.75,  283.75,
  283.85,    283.85,  283.85,  283.85,
  283.7,     283.7,   283.7,   283.7,
  283.35,    283.35,  283.35,  283.35,
  283,       283,     283,     283,
  282.65,    282.65,  282.65,  282.65,
  282.25,    282.25,  282.25,  282.25,
  282.05,    282.05,  282.05,  282.05,
  282.1,     282.1,   282.1,   282.1,
  281.95,    281.95,  281.95,  281.95,
  281.65,    281.65,  281.65,  281.65,
  281.4,     281.4,   281.4,   281.4,
  281,       281,     281,     281,
  280.55,    280.55,  280.55,  280.55,
  280.25,    280.25,  280.25,  280.25,
  280.3,     280.3,   280.3,   280.3,
  280.65,    280.65,  280.65,  280.65,
  281.3,     281.3,   281.3,   281.3,
  282.25,    282.25,  282.25,  282.25,
  283,       283,     283,     283,
  283.45,    283.45,  283.45,  283.45,
  284.1,     284.1,   284.1,   284.1,
  284.8,     284.8,   284.8,   284.8,
  285.1,     285.1,   285.1,   285.1,
  285.15,    285.15,  285.15,  285.15,
  285.35,    285.35,  285.35,  285.35,
  285.7,     285.7,   285.7,   285.7,
  285.9,     285.9,   285.9,   285.9,
  286.2,     286.2,   286.2,   286.2,
  286.4,     286.4,   286.4,   286.4,
  286.5,     286.5,   286.5,   286.5,
  286.5,     286.5,   286.5,   286.5,
  286.4,     286.4,   286.4,   286.4,
  286.4,     286.4,   286.4,   286.4,
  286.25,    286.25,  286.25,  286.25,
  286,       286,     286,     286,
  285.75,    285.75,  285.75,  285.75,
  285.65,    285.65,  285.65,  285.65,
  285.7,     285.7,   285.7,   285.7,
  285.7,     285.7,   285.7,   285.7,
  285.4,     285.4,   285.4,   285.4,
  284.85,    284.85,  284.85,  284.85,
  284.5,     284.5,   284.5,   284.5,
  284.5,     284.5,   284.5,   284.5,
  284.55,    284.55,  284.55,  284.55,
  284.55,    284.55,  284.55,  284.55,
  284.55,    284.55,  284.55,  284.55,
  284.3,     284.3,   284.3,   284.3,
  284,       284,     284,     284,
  284,       284,     284,     284,
  284,       284,     284,     284,
  283.65,    283.65,  283.65,  283.65,
  282.65,    282.65,  282.65,  282.65,
  280.95,    280.95,  280.95,  280.95,
  279.8,     279.8,   279.8,   279.8,
  279.65,    279.65,  279.65,  279.65,
  279.35,    279.35,  279.35,  279.35,
  278.95,    278.95,  278.95,  278.95,
  278.8,     278.8,   278.8,   278.8,
  278.7,     278.7,   278.7,   278.7,
  278.85,    278.85,  278.85,  278.85,
  279.2,     279.2,   279.2,   279.2,
  279.45,    279.45,  279.45,  279.45,
  279.65,    279.65,  279.65,  279.65,
  279.8,     279.8,   279.8,   279.8,
  279.85,    279.85,  279.85,  279.85,
  279.95,    279.95,  279.95,  279.95,
  280.15,    280.15,  280.15,  280.15,
  280.4,     280.4,   280.4,   280.4,
  280.6,     280.6,   280.6,   280.6,
  280.75,    280.75,  280.75,  280.75,
  280.9,     280.9,   280.9,   280.9,
  281,       281,     281,     281,
  280.95,    280.95,  280.95,  280.95,
  281,       281,     281,     281,
  281,       281,     281,     281,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.65,    280.65,  280.65,  280.65,
  280.65,    280.65,  280.65,  280.65,
  280.8,     280.8,   280.8,   280.8,
  280.65,    280.65,  280.65,  280.65,
  280.3,     280.3,   280.3,   280.3,
  280.15,    280.15,  280.15,  280.15,
  280.1,     280.1,   280.1,   280.1,
  280.05,    280.05,  280.05,  280.05,
  280,       280,     280,     280,
  279.95,    279.95,  279.95,  279.95,
  279.9,     279.9,   279.9,   279.9,
  279.85,    279.85,  279.85,  279.85,
  279.8,     279.8,   279.8,   279.8,
  279.6,     279.6,   279.6,   279.6,
  279.25,    279.25,  279.25,  279.25,
  279.05,    279.05,  279.05,  279.05,
  279.05,    279.05,  279.05,  279.05,
  278.9,     278.9,   278.9,   278.9,
  278.75,    278.75,  278.75,  278.75,
  278.55,    278.55,  278.55,  278.55,
  278.25,    278.25,  278.25,  278.25,
  278.25,    278.25,  278.25,  278.25,
  278.2,     278.2,   278.2,   278.2,
  277.9,     277.9,   277.9,   277.9,
  277.75,    277.75,  277.75,  277.75,
  277.65,    277.65,  277.65,  277.65,
  277.5,     277.5,   277.5,   277.5,
  277.65,    277.65,  277.65,  277.65,
  278.1,     278.1,   278.1,   278.1,
  278.4,     278.4,   278.4,   278.4,
  278.5,     278.5,   278.5,   278.5,
  278.65,    278.65,  278.65,  278.65,
  278.8,     278.8,   278.8,   278.8,
  278.95,    278.95,  278.95,  278.95,
  279.15,    279.15,  279.15,  279.15,
  279.35,    279.35,  279.35,  279.35,
  279.4,     279.4,   279.4,   279.4,
  279.75,    279.75,  279.75,  279.75,
  280.45,    280.45,  280.45,  280.45,
  280.9,     280.9,   280.9,   280.9,
  281.15,    281.15,  281.15,  281.15,
  281.15,    281.15,  281.15,  281.15,
  280.55,    280.55,  280.55,  280.55,
  280.3,     280.3,   280.3,   280.3,
  280.65,    280.65,  280.65,  280.65,
  281.05,    281.05,  281.05,  281.05,
  281.35,    281.35,  281.35,  281.35,
  281.2,     281.2,   281.2,   281.2,
  281.15,    281.15,  281.15,  281.15,
  281.3,     281.3,   281.3,   281.3,
  281.4,     281.4,   281.4,   281.4,
  281.4,     281.4,   281.4,   281.4,
  281.2,     281.2,   281.2,   281.2,
  281,       281,     281,     281,
  280.9,     280.9,   280.9,   280.9,
  280.7,     280.7,   280.7,   280.7,
  280.35,    280.35,  280.35,  280.35,
  280.1,     280.1,   280.1,   280.1,
  279.9,     279.9,   279.9,   279.9,
  279.8,     279.8,   279.8,   279.8,
  279.9,     279.9,   279.9,   279.9,
  279.9,     279.9,   279.9,   279.9,
  279.85,    279.85,  279.85,  279.85,
  279.85,    279.85,  279.85,  279.85,
  279.9,     279.9,   279.9,   279.9,
  279.7,     279.7,   279.7,   279.7,
  279.5,     279.5,   279.5,   279.5,
  279.65,    279.65,  279.65,  279.65,
  279.75,    279.75,  279.75,  279.75,
  279.55,    279.55,  279.55,  279.55,
  279.15,    279.15,  279.15,  279.15,
  278.7,     278.7,   278.7,   278.7,
  278.35,    278.35,  278.35,  278.35,
  278.2,     278.2,   278.2,   278.2,
  278,       278,     278,     278,
  277.75,    277.75,  277.75,  277.75,
  277.6,     277.6,   277.6,   277.6,
  277.55,    277.55,  277.55,  277.55,
  277.6,     277.6,   277.6,   277.6,
  277.6,     277.6,   277.6,   277.6,
  277.8,     277.8,   277.8,   277.8,
  278.5,     278.5,   278.5,   278.5,
  279.3,     279.3,   279.3,   279.3,
  280.15,    280.15,  280.15,  280.15,
  281.2,     281.2,   281.2,   281.2,
  282.15,    282.15,  282.15,  282.15,
  282.65,    282.65,  282.65,  282.65,
  282.95,    282.95,  282.95,  282.95,
  283.45,    283.45,  283.45,  283.45,
  284.15,    284.15,  284.15,  284.15,
  284.65,    284.65,  284.65,  284.65,
  284.95,    284.95,  284.95,  284.95,
  285.15,    285.15,  285.15,  285.15,
  285.15,    285.15,  285.15,  285.15,
  285.25,    285.25,  285.25,  285.25,
  285.6,     285.6,   285.6,   285.6,
  285.7,     285.7,   285.7,   285.7,
  285.55,    285.55,  285.55,  285.55,
  285.6,     285.6,   285.6,   285.6,
  285.5,     285.5,   285.5,   285.5,
  285.15,    285.15,  285.15,  285.15,
  284.7,     284.7,   284.7,   284.7,
  284.1,     284.1,   284.1,   284.1,
  283.35,    283.35,  283.35,  283.35,
  282.45,    282.45,  282.45,  282.45,
  281.5,     281.5,   281.5,   281.5,
  280.65,    280.65,  280.65,  280.65,
  280,       280,     280,     280,
  279.45,    279.45,  279.45,  279.45,
  279,       279,     279,     279,
  278.65,    278.65,  278.65,  278.65,
  278.3,     278.3,   278.3,   278.3,
  278.05,    278.05,  278.05,  278.05,
  277.8,     277.8,   277.8,   277.8,
  277.4,     277.4,   277.4,   277.4,
  276.9,     276.9,   276.9,   276.9,
  276.45,    276.45,  276.45,  276.45,
  276.2,     276.2,   276.2,   276.2,
  275.95,    275.95,  275.95,  275.95,
  275.65,    275.65,  275.65,  275.65,
  275.15,    275.15,  275.15,  275.15,
  274.1,     274.1,   274.1,   274.1,
  273.25,    273.25,  273.25,  273.25,
  273.3,     273.3,   273.3,   273.3,
  273.65,    273.65,  273.65,  273.65,
  273.55,    273.55,  273.55,  273.55,
  273.05,    273.05,  273.05,  273.05,
  273,       273,     273,     273,
  273.55,    273.55,  273.55,  273.55,
  274.35,    274.35,  274.35,  274.35,
  275.7,     275.7,   275.7,   275.7,
  277.6,     277.6,   277.6,   277.6,
  279.85,    279.85,  279.85,  279.85,
  281.65,    281.65,  281.65,  281.65,
  282.6,     282.6,   282.6,   282.6,
  283.25,    283.25,  283.25,  283.25,
  283.95,    283.95,  283.95,  283.95,
  284.55,    284.55,  284.55,  284.55,
  284.95,    284.95,  284.95,  284.95,
  285.45,    285.45,  285.45,  285.45,
  285.85,    285.85,  285.85,  285.85,
  286.15,    286.15,  286.15,  286.15,
  286.45,    286.45,  286.45,  286.45,
  286.7,     286.7,   286.7,   286.7,
  286.85,    286.85,  286.85,  286.85,
  287,       287,     287,     287,
  287.1,     287.1,   287.1,   287.1,
  287,       287,     287,     287,
  286.8,     286.8,   286.8,   286.8,
  286.5,     286.5,   286.5,   286.5,
  286.05,    286.05,  286.05,  286.05,
  285.35,    285.35,  285.35,  285.35,
  284.4,     284.4,   284.4,   284.4,
  283.55,    283.55,  283.55,  283.55,
  282.9,     282.9,   282.9,   282.9,
  282.45,    282.45,  282.45,  282.45,
  282.35,    282.35,  282.35,  282.35,
  282,       282,     282,     282,
  281.2,     281.2,   281.2,   281.2,
  280.65,    280.65,  280.65,  280.65,
  280.45,    280.45,  280.45,  280.45,
  280,       280,     280,     280,
  279.15,    279.15,  279.15,  279.15,
  278.8,     278.8,   278.8,   278.8,
  278.75,    278.75,  278.75,  278.75,
  278.25,    278.25,  278.25,  278.25,
  277.75,    277.75,  277.75,  277.75,
  277.55,    277.55,  277.55,  277.55,
  277.55,    277.55,  277.55,  277.55,
  277.9,     277.9,   277.9,   277.9,
  278.05,    278.05,  278.05,  278.05,
  277.7,     277.7,   277.7,   277.7,
  277.65,    277.65,  277.65,  277.65,
  277.55,    277.55,  277.55,  277.55,
  277.3,     277.3,   277.3,   277.3,
  277.5,     277.5,   277.5,   277.5,
  277.6,     277.6,   277.6,   277.6,
  277.65,    277.65,  277.65,  277.65,
  278.7,     278.7,   278.7,   278.7,
  280.5,     280.5,   280.5,   280.5,
  282.25,    282.25,  282.25,  282.25,
  283.7,     283.7,   283.7,   283.7,
  284.75,    284.75,  284.75,  284.75,
  285.5,     285.5,   285.5,   285.5,
  286.15,    286.15,  286.15,  286.15,
  286.7,     286.7,   286.7,   286.7,
  287.1,     287.1,   287.1,   287.1,
  287.5,     287.5,   287.5,   287.5,
  288.05,    288.05,  288.05,  288.05,
  288.45,    288.45,  288.45,  288.45,
  288.8,     288.8,   288.8,   288.8,
  289.1,     289.1,   289.1,   289.1,
  289.1,     289.1,   289.1,   289.1,
  289.1,     289.1,   289.1,   289.1,
  289.1,     289.1,   289.1,   289.1,
  288.95,    288.95,  288.95,  288.95,
  288.6,     288.6,   288.6,   288.6,
  288.1,     288.1,   288.1,   288.1,
  287.5,     287.5,   287.5,   287.5,
  286.7,     286.7,   286.7,   286.7,
  285.6,     285.6,   285.6,   285.6,
  284.5,     284.5,   284.5,   284.5,
  283.55,    283.55,  283.55,  283.55,
  282.55,    282.55,  282.55,  282.55,
  281.7,     281.7,   281.7,   281.7,
  281,       281,     281,     281,
  280.4,     280.4,   280.4,   280.4,
  280.25,    280.25,  280.25,  280.25,
  280.05,    280.05,  280.05,  280.05,
  279.45,    279.45,  279.45,  279.45,
  278.95,    278.95,  278.95,  278.95,
  278.6,     278.6,   278.6,   278.6,
  278.55,    278.55,  278.55,  278.55,
  278.55,    278.55,  278.55,  278.55,
  278.1,     278.1,   278.1,   278.1,
  277.75,    277.75,  277.75,  277.75,
  277.5,     277.5,   277.5,   277.5,
  277,       277,     277,     277,
  276.65,    276.65,  276.65,  276.65,
  276.2,     276.2,   276.2,   276.2,
  275.6,     275.6,   275.6,   275.6,
  275,       275,     275,     275,
  274.6,     274.6,   274.6,   274.6,
  274.75,    274.75,  274.75,  274.75,
  275.15,    275.15,  275.15,  275.15,
  275.85,    275.85,  275.85,  275.85,
  277.05,    277.05,  277.05,  277.05,
  278.35,    278.35,  278.35,  278.35,
  279.6,     279.6,   279.6,   279.6,
  280.9,     280.9,   280.9,   280.9,
  282.15,    282.15,  282.15,  282.15,
  283,       283,     283,     283,
  283.65,    283.65,  283.65,  283.65,
  284.15,    284.15,  284.15,  284.15,
  284.5,     284.5,   284.5,   284.5,
  284.9,     284.9,   284.9,   284.9,
  285.4,     285.4,   285.4,   285.4,
  285.85,    285.85,  285.85,  285.85,
  285.95,    285.95,  285.95,  285.95,
  286,       286,     286,     286,
  286.05,    286.05,  286.05,  286.05,
  286.05,    286.05,  286.05,  286.05,
  286,       286,     286,     286,
  285.95,    285.95,  285.95,  285.95,
  285.9,     285.9,   285.9,   285.9,
  285.8,     285.8,   285.8,   285.8,
  285.25,    285.25,  285.25,  285.25,
  284.65,    284.65,  284.65,  284.65,
  284.55,    284.55,  284.55,  284.55,
  284.5,     284.5,   284.5,   284.5,
  284.15,    284.15,  284.15,  284.15,
  283.45,    283.45,  283.45,  283.45,
  282.8,     282.8,   282.8,   282.8,
  282.4,     282.4,   282.4,   282.4,
  281.95,    281.95,  281.95,  281.95,
  280.8,     280.8,   280.8,   280.8,
  279.75,    279.75,  279.75,  279.75,
  279.75,    279.75,  279.75,  279.75,
  279.85,    279.85,  279.85,  279.85,
  279.9,     279.9,   279.9,   279.9,
  280.2,     280.2,   280.2,   280.2,
  280.4,     280.4,   280.4,   280.4,
  280.6,     280.6,   280.6,   280.6,
  280.9,     280.9,   280.9,   280.9,
  281.2,     281.2,   281.2,   281.2,
  281.4,     281.4,   281.4,   281.4,
  281.55,    281.55,  281.55,  281.55,
  281.6,     281.6,   281.6,   281.6,
  281.5,     281.5,   281.5,   281.5,
  281.55,    281.55,  281.55,  281.55,
  281.5,     281.5,   281.5,   281.5,
  281.1,     281.1,   281.1,   281.1,
  280.85,    280.85,  280.85,  280.85,
  281.05,    281.05,  281.05,  281.05,
  281.3,     281.3,   281.3,   281.3,
  281.7,     281.7,   281.7,   281.7,
  282.55,    282.55,  282.55,  282.55,
  283.25,    283.25,  283.25,  283.25,
  283.4,     283.4,   283.4,   283.4,
  283.35,    283.35,  283.35,  283.35,
  283.35,    283.35,  283.35,  283.35,
  283.6,     283.6,   283.6,   283.6,
  283.6,     283.6,   283.6,   283.6,
  283.1,     283.1,   283.1,   283.1,
  282.65,    282.65,  282.65,  282.65,
  282.3,     282.3,   282.3,   282.3,
  282.35,    282.35,  282.35,  282.35,
  282.85,    282.85,  282.85,  282.85,
  283.1,     283.1,   283.1,   283.1,
  282.9,     282.9,   282.9,   282.9,
  282.75,    282.75,  282.75,  282.75,
  282.55,    282.55,  282.55,  282.55,
  282.15,    282.15,  282.15,  282.15,
  281.9,     281.9,   281.9,   281.9,
  281.7,     281.7,   281.7,   281.7,
  281.35,    281.35,  281.35,  281.35,
  280.2,     280.2,   280.2,   280.2,
  279.2,     279.2,   279.2,   279.2,
  278.95,    278.95,  278.95,  278.95,
  278.6,     278.6,   278.6,   278.6,
  278.25,    278.25,  278.25,  278.25,
  277.95,    277.95,  277.95,  277.95,
  277.7,     277.7,   277.7,   277.7,
  277.35,    277.35,  277.35,  277.35,
  277.1,     277.1,   277.1,   277.1,
  276.95,    276.95,  276.95,  276.95,
  276.95,    276.95,  276.95,  276.95,
  277.25,    277.25,  277.25,  277.25,
  277.9,     277.9,   277.9,   277.9,
  278.15,    278.15,  278.15,  278.15,
  277.8,     277.8,   277.8,   277.8,
  277.55,    277.55,  277.55,  277.55,
  277.45,    277.45,  277.45,  277.45,
  277.4,     277.4,   277.4,   277.4,
  277.05,    277.05,  277.05,  277.05,
  276.75,    276.75,  276.75,  276.75,
  276.8,     276.8,   276.8,   276.8,
  276.85,    276.85,  276.85,  276.85,
  276.9,     276.9,   276.9,   276.9,
  277.1,     277.1,   277.1,   277.1,
  277.4,     277.4,   277.4,   277.4,
  277.4,     277.4,   277.4,   277.4,
  277.2,     277.2,   277.2,   277.2,
  277.95,    277.95,  277.95,  277.95,
  279,       279,     279,     279,
  278.85,    278.85,  278.85,  278.85,
  278.3,     278.3,   278.3,   278.3,
  278.95,    278.95,  278.95,  278.95,
  279.75,    279.75,  279.75,  279.75,
  280.05,    280.05,  280.05,  280.05,
  279.65,    279.65,  279.65,  279.65,
  279.55,    279.55,  279.55,  279.55,
  280.15,    280.15,  280.15,  280.15,
  280.25,    280.25,  280.25,  280.25,
  280.35,    280.35,  280.35,  280.35,
  279.65,    279.65,  279.65,  279.65,
  279.25,    279.25,  279.25,  279.25,
  279.35,    279.35,  279.35,  279.35,
  279.25,    279.25,  279.25,  279.25,
  279.35,    279.35,  279.35,  279.35,
  279.1,     279.1,   279.1,   279.1,
  278.95,    278.95,  278.95,  278.95,
  278.6,     278.6,   278.6,   278.6,
  278.1,     278.1,   278.1,   278.1,
  277.95,    277.95,  277.95,  277.95,
  277.55,    277.55,  277.55,  277.55,
  277.3,     277.3,   277.3,   277.3,
  277.35,    277.35,  277.35,  277.35,
  277.15,    277.15,  277.15,  277.15,
  276.7,     276.7,   276.7,   276.7,
  276.25,    276.25,  276.25,  276.25,
  276,       276,     276,     276,
  276.05,    276.05,  276.05,  276.05,
  276.35,    276.35,  276.35,  276.35,
  276.75,    276.75,  276.75,  276.75,
  277.05,    277.05,  277.05,  277.05,
  277.25,    277.25,  277.25,  277.25,
  277.4,     277.4,   277.4,   277.4,
  277.6,     277.6,   277.6,   277.6,
  277.8,     277.8,   277.8,   277.8,
  277.95,    277.95,  277.95,  277.95,
  278,       278,     278,     278,
  277.8,     277.8,   277.8,   277.8,
  277.8,     277.8,   277.8,   277.8,
  278.3,     278.3,   278.3,   278.3,
  279.05,    279.05,  279.05,  279.05,
  279.85,    279.85,  279.85,  279.85,
  280.65,    280.65,  280.65,  280.65,
  281.15,    281.15,  281.15,  281.15,
  281.3,     281.3,   281.3,   281.3,
  281.45,    281.45,  281.45,  281.45,
  281.6,     281.6,   281.6,   281.6,
  281.65,    281.65,  281.65,  281.65,
  281.6,     281.6,   281.6,   281.6,
  281.5,     281.5,   281.5,   281.5,
  281.5,     281.5,   281.5,   281.5,
  281.55,    281.55,  281.55,  281.55,
  281.55,    281.55,  281.55,  281.55,
  281.55,    281.55,  281.55,  281.55,
  281.6,     281.6,   281.6,   281.6,
  281.65,    281.65,  281.65,  281.65,
  281.65,    281.65,  281.65,  281.65,
  281.75,    281.75,  281.75,  281.75,
  281.9,     281.9,   281.9,   281.9,
  281.95,    281.95,  281.95,  281.95,
  282,       282,     282,     282,
  282.1,     282.1,   282.1,   282.1,
  282.2,     282.2,   282.2,   282.2,
  282.45,    282.45,  282.45,  282.45,
  282.9,     282.9,   282.9,   282.9,
  283.3,     283.3,   283.3,   283.3,
  283.5,     283.5,   283.5,   283.5,
  283.55,    283.55,  283.55,  283.55,
  283.5,     283.5,   283.5,   283.5,
  283.5,     283.5,   283.5,   283.5,
  283.65,    283.65,  283.65,  283.65,
  283.65,    283.65,  283.65,  283.65,
  283.35,    283.35,  283.35,  283.35,
  283,       283,     283,     283,
  282.05,    282.05,  282.05,  282.05,
  280.6,     280.6,   280.6,   280.6,
  279.8,     279.8,   279.8,   279.8,
  279.25,    279.25,  279.25,  279.25,
  278.5,     278.5,   278.5,   278.5,
  278.05,    278.05,  278.05,  278.05,
  277.85,    277.85,  277.85,  277.85,
  277.65,    277.65,  277.65,  277.65,
  277.5,     277.5,   277.5,   277.5,
  277.4,     277.4,   277.4,   277.4,
  277.3,     277.3,   277.3,   277.3,
  277.05,    277.05,  277.05,  277.05,
  276.55,    276.55,  276.55,  276.55,
  276.1,     276.1,   276.1,   276.1,
  275.75,    275.75,  275.75,  275.75,
  275.45,    275.45,  275.45,  275.45,
  275.25,    275.25,  275.25,  275.25,
  275.2,     275.2,   275.2,   275.2,
  275.85,    275.85,  275.85,  275.85,
  277.15,    277.15,  277.15,  277.15,
  278.2,     278.2,   278.2,   278.2,
  278.8,     278.8,   278.8,   278.8,
  279.3,     279.3,   279.3,   279.3,
  279.65,    279.65,  279.65,  279.65,
  279.95,    279.95,  279.95,  279.95,
  280.35,    280.35,  280.35,  280.35,
  280.7,     280.7,   280.7,   280.7,
  280.95,    280.95,  280.95,  280.95,
  281.1,     281.1,   281.1,   281.1,
  281.2,     281.2,   281.2,   281.2,
  281.2,     281.2,   281.2,   281.2,
  281.15,    281.15,  281.15,  281.15,
  281.2,     281.2,   281.2,   281.2,
  281.2,     281.2,   281.2,   281.2,
  281.15,    281.15,  281.15,  281.15,
  281.1,     281.1,   281.1,   281.1,
  281,       281,     281,     281,
  280.9,     280.9,   280.9,   280.9,
  280.65,    280.65,  280.65,  280.65,
  279.9,     279.9,   279.9,   279.9,
  279.2,     279.2,   279.2,   279.2,
  278.85,    278.85,  278.85,  278.85,
  278.2,     278.2,   278.2,   278.2,
  277.45,    277.45,  277.45,  277.45,
  276.7,     276.7,   276.7,   276.7,
  275.95,    275.95,  275.95,  275.95,
  275.4,     275.4,   275.4,   275.4,
  275.05,    275.05,  275.05,  275.05,
  274.7,     274.7,   274.7,   274.7,
  274.1,     274.1,   274.1,   274.1,
  273.6,     273.6,   273.6,   273.6,
  273.4,     273.4,   273.4,   273.4,
  273.4,     273.4,   273.4,   273.4,
  273.15,    273.15,  273.15,  273.15,
  272.65,    272.65,  272.65,  272.65,
  272.5,     272.5,   272.5,   272.5,
  272.45,    272.45,  272.45,  272.45,
  272,       272,     272,     272,
  271.55,    271.55,  271.55,  271.55,
  271.6,     271.6,   271.6,   271.6,
  271.2,     271.2,   271.2,   271.2,
  270.55,    270.55,  270.55,  270.55,
  270.75,    270.75,  270.75,  270.75,
  271.4,     271.4,   271.4,   271.4,
  271.9,     271.9,   271.9,   271.9,
  272.2,     272.2,   272.2,   272.2,
  272.9,     272.9,   272.9,   272.9,
  274.5,     274.5,   274.5,   274.5,
  276,       276,     276,     276,
  276.85,    276.85,  276.85,  276.85,
  277.6,     277.6,   277.6,   277.6,
  278.1,     278.1,   278.1,   278.1,
  278.55,    278.55,  278.55,  278.55,
  279.2,     279.2,   279.2,   279.2,
  279.65,    279.65,  279.65,  279.65,
  280.05,    280.05,  280.05,  280.05,
  280.65,    280.65,  280.65,  280.65,
  281.1,     281.1,   281.1,   281.1,
  281.35,    281.35,  281.35,  281.35,
  281.6,     281.6,   281.6,   281.6,
  281.95,    281.95,  281.95,  281.95,
  282.25,    282.25,  282.25,  282.25,
  282.4,     282.4,   282.4,   282.4,
  282.5,     282.5,   282.5,   282.5,
  282.5,     282.5,   282.5,   282.5,
  282.4,     282.4,   282.4,   282.4,
  282.3,     282.3,   282.3,   282.3,
  282.1,     282.1,   282.1,   282.1,
  281.7,     281.7,   281.7,   281.7,
  281.15,    281.15,  281.15,  281.15,
  280.45,    280.45,  280.45,  280.45,
  279.65,    279.65,  279.65,  279.65,
  278.85,    278.85,  278.85,  278.85,
  278.25,    278.25,  278.25,  278.25,
  277.8,     277.8,   277.8,   277.8,
  277.15,    277.15,  277.15,  277.15,
  276.8,     276.8,   276.8,   276.8,
  276.75,    276.75,  276.75,  276.75,
  276.7,     276.7,   276.7,   276.7,
  276.4,     276.4,   276.4,   276.4,
  275.8,     275.8,   275.8,   275.8,
  275.6,     275.6,   275.6,   275.6,
  275.55,    275.55,  275.55,  275.55,
  275.3,     275.3,   275.3,   275.3,
  275.25,    275.25,  275.25,  275.25,
  275.35,    275.35,  275.35,  275.35,
  275.15,    275.15,  275.15,  275.15,
  274.85,    274.85,  274.85,  274.85,
  274.55,    274.55,  274.55,  274.55,
  274.2,     274.2,   274.2,   274.2,
  274.05,    274.05,  274.05,  274.05,
  273.75,    273.75,  273.75,  273.75,
  273.7,     273.7,   273.7,   273.7,
  274.75,    274.75,  274.75,  274.75,
  276.3,     276.3,   276.3,   276.3,
  277.85,    277.85,  277.85,  277.85,
  279.3,     279.3,   279.3,   279.3,
  280.35,    280.35,  280.35,  280.35,
  281.25,    281.25,  281.25,  281.25,
  282.1,     282.1,   282.1,   282.1,
  282.7,     282.7,   282.7,   282.7,
  283.45,    283.45,  283.45,  283.45,
  284.15,    284.15,  284.15,  284.15,
  284.55,    284.55,  284.55,  284.55,
  285.1,     285.1,   285.1,   285.1,
  285.45,    285.45,  285.45,  285.45,
  285.7,     285.7,   285.7,   285.7,
  286.25,    286.25,  286.25,  286.25,
  286.7,     286.7,   286.7,   286.7,
  287,       287,     287,     287,
  287.2,     287.2,   287.2,   287.2,
  287.15,    287.15,  287.15,  287.15,
  286.85,    286.85,  286.85,  286.85,
  286.55,    286.55,  286.55,  286.55,
  286.35,    286.35,  286.35,  286.35,
  286,       286,     286,     286,
  285.35,    285.35,  285.35,  285.35,
  284.6,     284.6,   284.6,   284.6,
  283.8,     283.8,   283.8,   283.8,
  282.85,    282.85,  282.85,  282.85,
  282.05,    282.05,  282.05,  282.05,
  281.5,     281.5,   281.5,   281.5,
  281.1,     281.1,   281.1,   281.1,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.8,     280.8,   280.8,   280.8,
  280.9,     280.9,   280.9,   280.9,
  280.85,    280.85,  280.85,  280.85,
  280.55,    280.55,  280.55,  280.55,
  280.1,     280.1,   280.1,   280.1,
  279.65,    279.65,  279.65,  279.65,
  279.4,     279.4,   279.4,   279.4,
  279.25,    279.25,  279.25,  279.25,
  279.1,     279.1,   279.1,   279.1,
  279,       279,     279,     279,
  278.85,    278.85,  278.85,  278.85,
  278.6,     278.6,   278.6,   278.6,
  278.4,     278.4,   278.4,   278.4,
  278.5,     278.5,   278.5,   278.5,
  278.8,     278.8,   278.8,   278.8,
  279.35,    279.35,  279.35,  279.35,
  280.25,    280.25,  280.25,  280.25,
  281.3,     281.3,   281.3,   281.3,
  282.25,    282.25,  282.25,  282.25,
  282.95,    282.95,  282.95,  282.95,
  284,       284,     284,     284,
  285.2,     285.2,   285.2,   285.2,
  286.15,    286.15,  286.15,  286.15,
  286.85,    286.85,  286.85,  286.85,
  287.45,    287.45,  287.45,  287.45,
  288.15,    288.15,  288.15,  288.15,
  288.6,     288.6,   288.6,   288.6,
  288.9,     288.9,   288.9,   288.9,
  289.1,     289.1,   289.1,   289.1,
  289.4,     289.4,   289.4,   289.4,
  289.7,     289.7,   289.7,   289.7,
  289.7,     289.7,   289.7,   289.7,
  289.75,    289.75,  289.75,  289.75,
  289.95,    289.95,  289.95,  289.95,
  290.1,     290.1,   290.1,   290.1,
  290,       290,     290,     290,
  289.65,    289.65,  289.65,  289.65,
  289,       289,     289,     289,
  287.8,     287.8,   287.8,   287.8,
  286.35,    286.35,  286.35,  286.35,
  285.2,     285.2,   285.2,   285.2,
  284.35,    284.35,  284.35,  284.35,
  283.5,     283.5,   283.5,   283.5,
  283,       283,     283,     283,
  282.5,     282.5,   282.5,   282.5,
  281.6,     281.6,   281.6,   281.6,
  281,       281,     281,     281,
  280.35,    280.35,  280.35,  280.35,
  279.5,     279.5,   279.5,   279.5,
  278.95,    278.95,  278.95,  278.95,
  278.65,    278.65,  278.65,  278.65,
  278.35,    278.35,  278.35,  278.35,
  278.15,    278.15,  278.15,  278.15,
  278.05,    278.05,  278.05,  278.05,
  277.7,     277.7,   277.7,   277.7,
  277.2,     277.2,   277.2,   277.2,
  276.55,    276.55,  276.55,  276.55,
  275.95,    275.95,  275.95,  275.95,
  275.85,    275.85,  275.85,  275.85,
  275.6,     275.6,   275.6,   275.6,
  275.2,     275.2,   275.2,   275.2,
  275,       275,     275,     275,
  274.8,     274.8,   274.8,   274.8,
  274.85,    274.85,  274.85,  274.85,
  275.45,    275.45,  275.45,  275.45,
  276.65,    276.65,  276.65,  276.65,
  278.15,    278.15,  278.15,  278.15,
  279.55,    279.55,  279.55,  279.55,
  280.75,    280.75,  280.75,  280.75,
  282.35,    282.35,  282.35,  282.35,
  283.8,     283.8,   283.8,   283.8,
  284.75,    284.75,  284.75,  284.75,
  285.65,    285.65,  285.65,  285.65,
  286.3,     286.3,   286.3,   286.3,
  286.85,    286.85,  286.85,  286.85,
  287.4,     287.4,   287.4,   287.4,
  287.85,    287.85,  287.85,  287.85,
  288.2,     288.2,   288.2,   288.2,
  288.4,     288.4,   288.4,   288.4,
  288.55,    288.55,  288.55,  288.55,
  288.7,     288.7,   288.7,   288.7,
  288.7,     288.7,   288.7,   288.7,
  288.6,     288.6,   288.6,   288.6,
  288.4,     288.4,   288.4,   288.4,
  288,       288,     288,     288,
  287.5,     287.5,   287.5,   287.5,
  286.8,     286.8,   286.8,   286.8,
  285.8,     285.8,   285.8,   285.8,
  284.6,     284.6,   284.6,   284.6,
  283.5,     283.5,   283.5,   283.5,
  282.9,     282.9,   282.9,   282.9,
  282.35,    282.35,  282.35,  282.35,
  281.45,    281.45,  281.45,  281.45,
  280.75,    280.75,  280.75,  280.75,
  280.15,    280.15,  280.15,  280.15,
  279.5,     279.5,   279.5,   279.5,
  279.05,    279.05,  279.05,  279.05,
  278.6,     278.6,   278.6,   278.6,
  278.15,    278.15,  278.15,  278.15,
  277.8,     277.8,   277.8,   277.8,
  277.7,     277.7,   277.7,   277.7,
  277.75,    277.75,  277.75,  277.75,
  277.65,    277.65,  277.65,  277.65,
  277.5,     277.5,   277.5,   277.5,
  277.6,     277.6,   277.6,   277.6,
  278.1,     278.1,   278.1,   278.1,
  278.85,    278.85,  278.85,  278.85,
  279.45,    279.45,  279.45,  279.45,
  279.8,     279.8,   279.8,   279.8,
  280.05,    280.05,  280.05,  280.05,
  280.35,    280.35,  280.35,  280.35,
  280.8,     280.8,   280.8,   280.8,
  281.3,     281.3,   281.3,   281.3,
  281.85,    281.85,  281.85,  281.85,
  282.4,     282.4,   282.4,   282.4,
  282.5,     282.5,   282.5,   282.5,
  282,       282,     282,     282,
  281.7,     281.7,   281.7,   281.7,
  281.7,     281.7,   281.7,   281.7,
  280.95,    280.95,  280.95,  280.95,
  280.35,    280.35,  280.35,  280.35,
  280.4,     280.4,   280.4,   280.4,
  280.35,    280.35,  280.35,  280.35,
  280.35,    280.35,  280.35,  280.35,
  280.45,    280.45,  280.45,  280.45,
  280.3,     280.3,   280.3,   280.3,
  280.3,     280.3,   280.3,   280.3,
  280.7,     280.7,   280.7,   280.7,
  280.65,    280.65,  280.65,  280.65,
  280.4,     280.4,   280.4,   280.4,
  280.25,    280.25,  280.25,  280.25,
  280.2,     280.2,   280.2,   280.2,
  280.2,     280.2,   280.2,   280.2,
  280.1,     280.1,   280.1,   280.1,
  280,       280,     280,     280,
  279.9,     279.9,   279.9,   279.9,
  279.65,    279.65,  279.65,  279.65,
  279.35,    279.35,  279.35,  279.35,
  279.2,     279.2,   279.2,   279.2,
  279.15,    279.15,  279.15,  279.15,
  279,       279,     279,     279,
  278.7,     278.7,   278.7,   278.7,
  278.4,     278.4,   278.4,   278.4,
  278.4,     278.4,   278.4,   278.4,
  278.6,     278.6,   278.6,   278.6,
  278.55,    278.55,  278.55,  278.55,
  278.4,     278.4,   278.4,   278.4,
  278.45,    278.45,  278.45,  278.45,
  278.5,     278.5,   278.5,   278.5,
  278.1,     278.1,   278.1,   278.1,
  277.7,     277.7,   277.7,   277.7,
  277.55,    277.55,  277.55,  277.55,
  277.3,     277.3,   277.3,   277.3,
  277.05,    277.05,  277.05,  277.05,
  277,       277,     277,     277,
  277.2,     277.2,   277.2,   277.2,
  277.3,     277.3,   277.3,   277.3,
  277.45,    277.45,  277.45,  277.45,
  278,       278,     278,     278,
  278.65,    278.65,  278.65,  278.65,
  278.95,    278.95,  278.95,  278.95,
  278.95,    278.95,  278.95,  278.95,
  278.9,     278.9,   278.9,   278.9,
  278.95,    278.95,  278.95,  278.95,
  279.4,     279.4,   279.4,   279.4,
  279.6,     279.6,   279.6,   279.6,
  279.5,     279.5,   279.5,   279.5,
  280.25,    280.25,  280.25,  280.25,
  280.9,     280.9,   280.9,   280.9,
  280.9,     280.9,   280.9,   280.9,
  281.2,     281.2,   281.2,   281.2,
  281.5,     281.5,   281.5,   281.5,
  281.6,     281.6,   281.6,   281.6,
  281.45,    281.45,  281.45,  281.45,
  281.25,    281.25,  281.25,  281.25,
  281.25,    281.25,  281.25,  281.25,
  281,       281,     281,     281,
  280.7,     280.7,   280.7,   280.7,
  280.4,     280.4,   280.4,   280.4,
  280,       280,     280,     280,
  279.8,     279.8,   279.8,   279.8,
  279.6,     279.6,   279.6,   279.6,
  279.1,     279.1,   279.1,   279.1,
  278.25,    278.25,  278.25,  278.25,
  277.85,    277.85,  277.85,  277.85,
  277.9,     277.9,   277.9,   277.9,
  277.65,    277.65,  277.65,  277.65,
  277.3,     277.3,   277.3,   277.3,
  276.9,     276.9,   276.9,   276.9,
  276.55,    276.55,  276.55,  276.55,
  276.25,    276.25,  276.25,  276.25,
  275.85,    275.85,  275.85,  275.85,
  275.4,     275.4,   275.4,   275.4,
  274.85,    274.85,  274.85,  274.85,
  274.2,     274.2,   274.2,   274.2,
  273.65,    273.65,  273.65,  273.65,
  273.45,    273.45,  273.45,  273.45,
  273.4,     273.4,   273.4,   273.4,
  273.25,    273.25,  273.25,  273.25,
  273.3,     273.3,   273.3,   273.3,
  273.55,    273.55,  273.55,  273.55,
  273.7,     273.7,   273.7,   273.7,
  273.6,     273.6,   273.6,   273.6,
  273.2,     273.2,   273.2,   273.2,
  272.65,    272.65,  272.65,  272.65,
  272.55,    272.55,  272.55,  272.55,
  272.9,     272.9,   272.9,   272.9,
  273.65,    273.65,  273.65,  273.65,
  275.25,    275.25,  275.25,  275.25,
  277.3,     277.3,   277.3,   277.3,
  278.85,    278.85,  278.85,  278.85,
  279.65,    279.65,  279.65,  279.65,
  279.95,    279.95,  279.95,  279.95,
  280.3,     280.3,   280.3,   280.3,
  280.65,    280.65,  280.65,  280.65,
  280.85,    280.85,  280.85,  280.85,
  281.3,     281.3,   281.3,   281.3,
  281.85,    281.85,  281.85,  281.85,
  282.35,    282.35,  282.35,  282.35,
  282.7,     282.7,   282.7,   282.7,
  282.95,    282.95,  282.95,  282.95,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  282.95,    282.95,  282.95,  282.95,
  282.35,    282.35,  282.35,  282.35,
  281.9,     281.9,   281.9,   281.9,
  281.55,    281.55,  281.55,  281.55,
  281.15,    281.15,  281.15,  281.15,
  280.85,    280.85,  280.85,  280.85,
  280.65,    280.65,  280.65,  280.65,
  280.5,     280.5,   280.5,   280.5,
  280.35,    280.35,  280.35,  280.35,
  280.15,    280.15,  280.15,  280.15,
  280,       280,     280,     280,
  279.9,     279.9,   279.9,   279.9,
  279.85,    279.85,  279.85,  279.85,
  279.8,     279.8,   279.8,   279.8,
  279.7,     279.7,   279.7,   279.7,
  279.6,     279.6,   279.6,   279.6,
  279.5,     279.5,   279.5,   279.5,
  279.4,     279.4,   279.4,   279.4,
  279.35,    279.35,  279.35,  279.35,
  279.35,    279.35,  279.35,  279.35,
  279.4,     279.4,   279.4,   279.4,
  279.5,     279.5,   279.5,   279.5,
  279.65,    279.65,  279.65,  279.65,
  279.8,     279.8,   279.8,   279.8,
  279.75,    279.75,  279.75,  279.75,
  279.6,     279.6,   279.6,   279.6,
  279.5,     279.5,   279.5,   279.5,
  279.45,    279.45,  279.45,  279.45,
  279.5,     279.5,   279.5,   279.5,
  279.55,    279.55,  279.55,  279.55,
  279.75,    279.75,  279.75,  279.75,
  280.25,    280.25,  280.25,  280.25,
  280.65,    280.65,  280.65,  280.65,
  280.9,     280.9,   280.9,   280.9,
  281.4,     281.4,   281.4,   281.4,
  282.25,    282.25,  282.25,  282.25,
  283.25,    283.25,  283.25,  283.25,
  284.05,    284.05,  284.05,  284.05,
  284.35,    284.35,  284.35,  284.35,
  284.3,     284.3,   284.3,   284.3,
  283.8,     283.8,   283.8,   283.8,
  283.05,    283.05,  283.05,  283.05,
  282.65,    282.65,  282.65,  282.65,
  282.8,     282.8,   282.8,   282.8,
  283.05,    283.05,  283.05,  283.05,
  282.75,    282.75,  282.75,  282.75,
  282.35,    282.35,  282.35,  282.35,
  282.2,     282.2,   282.2,   282.2,
  282.05,    282.05,  282.05,  282.05,
  282,       282,     282,     282,
  282.05,    282.05,  282.05,  282.05,
  281.95,    281.95,  281.95,  281.95,
  281.65,    281.65,  281.65,  281.65,
  281.2,     281.2,   281.2,   281.2,
  280.65,    280.65,  280.65,  280.65,
  280.1,     280.1,   280.1,   280.1,
  279.7,     279.7,   279.7,   279.7,
  279.55,    279.55,  279.55,  279.55,
  279.5,     279.5,   279.5,   279.5,
  279.4,     279.4,   279.4,   279.4,
  279.25,    279.25,  279.25,  279.25,
  279.1,     279.1,   279.1,   279.1,
  278.8,     278.8,   278.8,   278.8,
  278.6,     278.6,   278.6,   278.6,
  278.65,    278.65,  278.65,  278.65,
  278.65,    278.65,  278.65,  278.65,
  278.6,     278.6,   278.6,   278.6,
  278.55,    278.55,  278.55,  278.55,
  278.5,     278.5,   278.5,   278.5,
  278.4,     278.4,   278.4,   278.4,
  278.2,     278.2,   278.2,   278.2,
  277.9,     277.9,   277.9,   277.9,
  277.85,    277.85,  277.85,  277.85,
  277.7,     277.7,   277.7,   277.7,
  277.4,     277.4,   277.4,   277.4,
  277.25,    277.25,  277.25,  277.25,
  277.2,     277.2,   277.2,   277.2,
  277.15,    277.15,  277.15,  277.15,
  277.45,    277.45,  277.45,  277.45,
  278.05,    278.05,  278.05,  278.05,
  278.6,     278.6,   278.6,   278.6,
  279.1,     279.1,   279.1,   279.1,
  279.5,     279.5,   279.5,   279.5,
  279.85,    279.85,  279.85,  279.85,
  280,       280,     280,     280,
  280.25,    280.25,  280.25,  280.25,
  280.6,     280.6,   280.6,   280.6,
  280.8,     280.8,   280.8,   280.8,
  280.95,    280.95,  280.95,  280.95,
  281.1,     281.1,   281.1,   281.1,
  281.4,     281.4,   281.4,   281.4,
  281.6,     281.6,   281.6,   281.6,
  281.5,     281.5,   281.5,   281.5,
  281.45,    281.45,  281.45,  281.45,
  281.35,    281.35,  281.35,  281.35,
  281.15,    281.15,  281.15,  281.15,
  281.05,    281.05,  281.05,  281.05,
  280.7,     280.7,   280.7,   280.7,
  280.3,     280.3,   280.3,   280.3,
  280.15,    280.15,  280.15,  280.15,
  279.9,     279.9,   279.9,   279.9,
  279.7,     279.7,   279.7,   279.7,
  279.45,    279.45,  279.45,  279.45,
  278.85,    278.85,  278.85,  278.85,
  278.3,     278.3,   278.3,   278.3,
  278.05,    278.05,  278.05,  278.05,
  277.7,     277.7,   277.7,   277.7,
  277.3,     277.3,   277.3,   277.3,
  277,       277,     277,     277,
  276.85,    276.85,  276.85,  276.85,
  276.7,     276.7,   276.7,   276.7,
  276.45,    276.45,  276.45,  276.45,
  276.4,     276.4,   276.4,   276.4,
  276.35,    276.35,  276.35,  276.35,
  276.1,     276.1,   276.1,   276.1,
  276,       276,     276,     276,
  275.9,     275.9,   275.9,   275.9,
  275.8,     275.8,   275.8,   275.8,
  275.95,    275.95,  275.95,  275.95,
  276.2,     276.2,   276.2,   276.2,
  276.3,     276.3,   276.3,   276.3,
  276.2,     276.2,   276.2,   276.2,
  276.3,     276.3,   276.3,   276.3,
  276.35,    276.35,  276.35,  276.35,
  276.35,    276.35,  276.35,  276.35,
  276.55,    276.55,  276.55,  276.55,
  276.8,     276.8,   276.8,   276.8,
  277.2,     277.2,   277.2,   277.2,
  277.75,    277.75,  277.75,  277.75,
  278.35,    278.35,  278.35,  278.35,
  278.85,    278.85,  278.85,  278.85,
  279.25,    279.25,  279.25,  279.25,
  279.6,     279.6,   279.6,   279.6,
  279.85,    279.85,  279.85,  279.85,
  280.25,    280.25,  280.25,  280.25,
  280.9,     280.9,   280.9,   280.9,
  281.25,    281.25,  281.25,  281.25,
  281.5,     281.5,   281.5,   281.5,
  281.9,     281.9,   281.9,   281.9,
  281.95,    281.95,  281.95,  281.95,
  281.75,    281.75,  281.75,  281.75,
  281.7,     281.7,   281.7,   281.7,
  281.8,     281.8,   281.8,   281.8,
  282.05,    282.05,  282.05,  282.05,
  282.2,     282.2,   282.2,   282.2,
  282.2,     282.2,   282.2,   282.2,
  282.05,    282.05,  282.05,  282.05,
  281.7,     281.7,   281.7,   281.7,
  281.45,    281.45,  281.45,  281.45,
  281.2,     281.2,   281.2,   281.2,
  280.8,     280.8,   280.8,   280.8,
  280.35,    280.35,  280.35,  280.35,
  280.05,    280.05,  280.05,  280.05,
  279.8,     279.8,   279.8,   279.8,
  279.4,     279.4,   279.4,   279.4,
  279,       279,     279,     279,
  278.65,    278.65,  278.65,  278.65,
  278.2,     278.2,   278.2,   278.2,
  277.75,    277.75,  277.75,  277.75,
  277.25,    277.25,  277.25,  277.25,
  276.75,    276.75,  276.75,  276.75,
  276.35,    276.35,  276.35,  276.35,
  276,       276,     276,     276,
  275.6,     275.6,   275.6,   275.6,
  275.2,     275.2,   275.2,   275.2,
  275,       275,     275,     275,
  274.95,    274.95,  274.95,  274.95,
  274.85,    274.85,  274.85,  274.85,
  274.6,     274.6,   274.6,   274.6,
  274.25,    274.25,  274.25,  274.25,
  273.9,     273.9,   273.9,   273.9,
  273.65,    273.65,  273.65,  273.65,
  273.65,    273.65,  273.65,  273.65,
  273.85,    273.85,  273.85,  273.85,
  274.2,     274.2,   274.2,   274.2,
  275.4,     275.4,   275.4,   275.4,
  277.15,    277.15,  277.15,  277.15,
  278.8,     278.8,   278.8,   278.8,
  280.45,    280.45,  280.45,  280.45,
  281.65,    281.65,  281.65,  281.65,
  282.25,    282.25,  282.25,  282.25,
  282.7,     282.7,   282.7,   282.7,
  283.2,     283.2,   283.2,   283.2,
  283.6,     283.6,   283.6,   283.6,
  283.9,     283.9,   283.9,   283.9,
  284.25,    284.25,  284.25,  284.25,
  284.7,     284.7,   284.7,   284.7,
  285.15,    285.15,  285.15,  285.15,
  285.35,    285.35,  285.35,  285.35,
  285.5,     285.5,   285.5,   285.5,
  285.7,     285.7,   285.7,   285.7,
  285.8,     285.8,   285.8,   285.8,
  285.8,     285.8,   285.8,   285.8,
  285.5,     285.5,   285.5,   285.5,
  285.1,     285.1,   285.1,   285.1,
  284.6,     284.6,   284.6,   284.6,
  284.1,     284.1,   284.1,   284.1,
  283.65,    283.65,  283.65,  283.65,
  283,       283,     283,     283,
  282.2,     282.2,   282.2,   282.2,
  281.3,     281.3,   281.3,   281.3,
  280.5,     280.5,   280.5,   280.5,
  279.8,     279.8,   279.8,   279.8,
  279.1,     279.1,   279.1,   279.1,
  278.5,     278.5,   278.5,   278.5,
  278.15,    278.15,  278.15,  278.15,
  277.8,     277.8,   277.8,   277.8,
  277.1,     277.1,   277.1,   277.1,
  276.5,     276.5,   276.5,   276.5,
  276.15,    276.15,  276.15,  276.15,
  275.75,    275.75,  275.75,  275.75,
  275.35,    275.35,  275.35,  275.35,
  275.05,    275.05,  275.05,  275.05,
  274.7,     274.7,   274.7,   274.7,
  274.45,    274.45,  274.45,  274.45,
  274.35,    274.35,  274.35,  274.35,
  273.95,    273.95,  273.95,  273.95,
  273.5,     273.5,   273.5,   273.5,
  273,       273,     273,     273,
  272.75,    272.75,  272.75,  272.75,
  273.15,    273.15,  273.15,  273.15,
  273.4,     273.4,   273.4,   273.4,
  273.8,     273.8,   273.8,   273.8,
  274.95,    274.95,  274.95,  274.95,
  276.5,     276.5,   276.5,   276.5,
  277.9,     277.9,   277.9,   277.9,
  278.85,    278.85,  278.85,  278.85,
  279.35,    279.35,  279.35,  279.35,
  279.65,    279.65,  279.65,  279.65,
  279.85,    279.85,  279.85,  279.85,
  279.7,     279.7,   279.7,   279.7,
  279.95,    279.95,  279.95,  279.95,
  280.55,    280.55,  280.55,  280.55,
  280.75,    280.75,  280.75,  280.75,
  280.8,     280.8,   280.8,   280.8,
  280.8,     280.8,   280.8,   280.8,
  281.25,    281.25,  281.25,  281.25,
  281.9,     281.9,   281.9,   281.9,
  282.1,     282.1,   282.1,   282.1,
  282.45,    282.45,  282.45,  282.45,
  282.7,     282.7,   282.7,   282.7,
  282.75,    282.75,  282.75,  282.75,
  282.7,     282.7,   282.7,   282.7,
  282.6,     282.6,   282.6,   282.6,
  282.45,    282.45,  282.45,  282.45,
  281.9,     281.9,   281.9,   281.9,
  281.15,    281.15,  281.15,  281.15,
  280.25,    280.25,  280.25,  280.25,
  279.4,     279.4,   279.4,   279.4,
  278.8,     278.8,   278.8,   278.8,
  278.4,     278.4,   278.4,   278.4,
  278.35,    278.35,  278.35,  278.35,
  278.7,     278.7,   278.7,   278.7,
  279.05,    279.05,  279.05,  279.05,
  279.1,     279.1,   279.1,   279.1,
  278.95,    278.95,  278.95,  278.95,
  278.8,     278.8,   278.8,   278.8,
  278.7,     278.7,   278.7,   278.7,
  278.6,     278.6,   278.6,   278.6,
  278.45,    278.45,  278.45,  278.45,
  278.25,    278.25,  278.25,  278.25,
  278,       278,     278,     278,
  277.75,    277.75,  277.75,  277.75,
  277.55,    277.55,  277.55,  277.55,
  277.35,    277.35,  277.35,  277.35,
  277.2,     277.2,   277.2,   277.2,
  277.2,     277.2,   277.2,   277.2,
  277.3,     277.3,   277.3,   277.3,
  277.45,    277.45,  277.45,  277.45,
  277.65,    277.65,  277.65,  277.65,
  277.95,    277.95,  277.95,  277.95,
  278.3,     278.3,   278.3,   278.3,
  278.45,    278.45,  278.45,  278.45,
  278.45,    278.45,  278.45,  278.45,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.5,     278.5,   278.5,   278.5,
  278.55,    278.55,  278.55,  278.55,
  278.7,     278.7,   278.7,   278.7,
  278.95,    278.95,  278.95,  278.95,
  279,       279,     279,     279,
  279,       279,     279,     279,
  279,       279,     279,     279,
  279.2,     279.2,   279.2,   279.2,
  279.2,     279.2,   279.2,   279.2,
  278.95,    278.95,  278.95,  278.95,
  279.3,     279.3,   279.3,   279.3,
  279.7,     279.7,   279.7,   279.7,
  279.7,     279.7,   279.7,   279.7,
  279.65,    279.65,  279.65,  279.65,
  279.9,     279.9,   279.9,   279.9,
  279.95,    279.95,  279.95,  279.95,
  279.8,     279.8,   279.8,   279.8,
  279.75,    279.75,  279.75,  279.75,
  279.3,     279.3,   279.3,   279.3,
  278.65,    278.65,  278.65,  278.65,
  278.2,     278.2,   278.2,   278.2,
  277.8,     277.8,   277.8,   277.8,
  277.5,     277.5,   277.5,   277.5,
  277.4,     277.4,   277.4,   277.4,
  277.35,    277.35,  277.35,  277.35,
  277.15,    277.15,  277.15,  277.15,
  276.65,    276.65,  276.65,  276.65,
  276.15,    276.15,  276.15,  276.15,
  275.65,    275.65,  275.65,  275.65,
  275.1,     275.1,   275.1,   275.1,
  274.65,    274.65,  274.65,  274.65,
  274.25,    274.25,  274.25,  274.25,
  273.9,     273.9,   273.9,   273.9,
  273.65,    273.65,  273.65,  273.65,
  273.4,     273.4,   273.4,   273.4,
  273.05,    273.05,  273.05,  273.05,
  272.65,    272.65,  272.65,  272.65,
  272.25,    272.25,  272.25,  272.25,
  271.95,    271.95,  271.95,  271.95,
  271.8,     271.8,   271.8,   271.8,
  271.9,     271.9,   271.9,   271.9,
  272.55,    272.55,  272.55,  272.55,
  273.75,    273.75,  273.75,  273.75,
  275.15,    275.15,  275.15,  275.15,
  276.3,     276.3,   276.3,   276.3,
  277.2,     277.2,   277.2,   277.2,
  277.85,    277.85,  277.85,  277.85,
  278.3,     278.3,   278.3,   278.3,
  278.45,    278.45,  278.45,  278.45,
  278.6,     278.6,   278.6,   278.6,
  279.05,    279.05,  279.05,  279.05,
  279.25,    279.25,  279.25,  279.25,
  279.45,    279.45,  279.45,  279.45,
  279.95,    279.95,  279.95,  279.95,
  280.3,     280.3,   280.3,   280.3,
  280.4,     280.4,   280.4,   280.4,
  280.3,     280.3,   280.3,   280.3,
  280.25,    280.25,  280.25,  280.25,
  280.5,     280.5,   280.5,   280.5,
  280.55,    280.55,  280.55,  280.55,
  280.3,     280.3,   280.3,   280.3,
  280.25,    280.25,  280.25,  280.25,
  280.1,     280.1,   280.1,   280.1,
  279.9,     279.9,   279.9,   279.9,
  279.75,    279.75,  279.75,  279.75,
  279.15,    279.15,  279.15,  279.15,
  278.45,    278.45,  278.45,  278.45,
  277.9,     277.9,   277.9,   277.9,
  277.25,    277.25,  277.25,  277.25,
  276.55,    276.55,  276.55,  276.55,
  276,       276,     276,     276,
  275.5,     275.5,   275.5,   275.5,
  275,       275,     275,     275,
  274.55,    274.55,  274.55,  274.55,
  274.2,     274.2,   274.2,   274.2,
  273.95,    273.95,  273.95,  273.95,
  273.6,     273.6,   273.6,   273.6,
  273.25,    273.25,  273.25,  273.25,
  273.1,     273.1,   273.1,   273.1,
  273,       273,     273,     273,
  272.95,    272.95,  272.95,  272.95,
  273,       273,     273,     273,
  272.9,     272.9,   272.9,   272.9,
  272.6,     272.6,   272.6,   272.6,
  272.5,     272.5,   272.5,   272.5,
  272.6,     272.6,   272.6,   272.6,
  272.6,     272.6,   272.6,   272.6,
  272.45,    272.45,  272.45,  272.45,
  272.35,    272.35,  272.35,  272.35,
  272.8,     272.8,   272.8,   272.8,
  274.15,    274.15,  274.15,  274.15,
  275.75,    275.75,  275.75,  275.75,
  277.05,    277.05,  277.05,  277.05,
  278,       278,     278,     278,
  278.7,     278.7,   278.7,   278.7,
  279.25,    279.25,  279.25,  279.25,
  279.85,    279.85,  279.85,  279.85,
  280.35,    280.35,  280.35,  280.35,
  280.55,    280.55,  280.55,  280.55,
  280.95,    280.95,  280.95,  280.95,
  281.55,    281.55,  281.55,  281.55,
  281.8,     281.8,   281.8,   281.8,
  281.9,     281.9,   281.9,   281.9,
  282.15,    282.15,  282.15,  282.15,
  282.25,    282.25,  282.25,  282.25,
  282.35,    282.35,  282.35,  282.35,
  282.5,     282.5,   282.5,   282.5,
  282.5,     282.5,   282.5,   282.5,
  282.4,     282.4,   282.4,   282.4,
  282.25,    282.25,  282.25,  282.25,
  282,       282,     282,     282,
  281.65,    281.65,  281.65,  281.65,
  281.2,     281.2,   281.2,   281.2,
  280.65,    280.65,  280.65,  280.65,
  279.9,     279.9,   279.9,   279.9,
  279.15,    279.15,  279.15,  279.15,
  278.7,     278.7,   278.7,   278.7,
  278.5,     278.5,   278.5,   278.5,
  278.45,    278.45,  278.45,  278.45,
  278.25,    278.25,  278.25,  278.25,
  277.9,     277.9,   277.9,   277.9,
  277.65,    277.65,  277.65,  277.65,
  277.45,    277.45,  277.45,  277.45,
  277.3,     277.3,   277.3,   277.3,
  277.35,    277.35,  277.35,  277.35,
  277.55,    277.55,  277.55,  277.55,
  277.65,    277.65,  277.65,  277.65,
  277.5,     277.5,   277.5,   277.5,
  277.1,     277.1,   277.1,   277.1,
  276.45,    276.45,  276.45,  276.45,
  275.8,     275.8,   275.8,   275.8,
  275.35,    275.35,  275.35,  275.35,
  275.1,     275.1,   275.1,   275.1,
  275.05,    275.05,  275.05,  275.05,
  275,       275,     275,     275,
  274.75,    274.75,  274.75,  274.75,
  274.45,    274.45,  274.45,  274.45,
  274.6,     274.6,   274.6,   274.6,
  275.5,     275.5,   275.5,   275.5,
  276.6,     276.6,   276.6,   276.6,
  277.85,    277.85,  277.85,  277.85,
  279.05,    279.05,  279.05,  279.05,
  279.15,    279.15,  279.15,  279.15,
  278.6,     278.6,   278.6,   278.6,
  278.85,    278.85,  278.85,  278.85,
  279.9,     279.9,   279.9,   279.9,
  280.6,     280.6,   280.6,   280.6,
  280.8,     280.8,   280.8,   280.8,
  280.85,    280.85,  280.85,  280.85,
  280.8,     280.8,   280.8,   280.8,
  280.8,     280.8,   280.8,   280.8,
  281.2,     281.2,   281.2,   281.2,
  281.5,     281.5,   281.5,   281.5,
  281.45,    281.45,  281.45,  281.45,
  281.85,    281.85,  281.85,  281.85,
  282.3,     282.3,   282.3,   282.3,
  282.05,    282.05,  282.05,  282.05,
  281.35,    281.35,  281.35,  281.35,
  280.95,    280.95,  280.95,  280.95,
  280.9,     280.9,   280.9,   280.9,
  280.45,    280.45,  280.45,  280.45,
  280,       280,     280,     280,
  279.8,     279.8,   279.8,   279.8,
  279.35,    279.35,  279.35,  279.35,
  278.75,    278.75,  278.75,  278.75,
  278.15,    278.15,  278.15,  278.15,
  277.5,     277.5,   277.5,   277.5,
  277,       277,     277,     277,
  276.85,    276.85,  276.85,  276.85,
  276.65,    276.65,  276.65,  276.65,
  276.15,    276.15,  276.15,  276.15,
  275.75,    275.75,  275.75,  275.75,
  275.4,     275.4,   275.4,   275.4,
  274.7,     274.7,   274.7,   274.7,
  274,       274,     274,     274,
  273.6,     273.6,   273.6,   273.6,
  272.7,     272.7,   272.7,   272.7,
  272.9,     272.9,   272.9,   272.9,
  273.8,     273.8,   273.8,   273.8,
  273.45,    273.45,  273.45,  273.45,
  272.75,    272.75,  272.75,  272.75,
  272.4,     272.4,   272.4,   272.4,
  272.45,    272.45,  272.45,  272.45,
  272.35,    272.35,  272.35,  272.35,
  271.8,     271.8,   271.8,   271.8,
  271.6,     271.6,   271.6,   271.6,
  272.6,     272.6,   272.6,   272.6,
  274.5,     274.5,   274.5,   274.5,
  276.65,    276.65,  276.65,  276.65,
  278.2,     278.2,   278.2,   278.2,
  279.1,     279.1,   279.1,   279.1,
  279.85,    279.85,  279.85,  279.85,
  280.45,    280.45,  280.45,  280.45,
  281.05,    281.05,  281.05,  281.05,
  281.65,    281.65,  281.65,  281.65,
  282.15,    282.15,  282.15,  282.15,
  282.7,     282.7,   282.7,   282.7,
  283.1,     283.1,   283.1,   283.1,
  283.45,    283.45,  283.45,  283.45,
  283.8,     283.8,   283.8,   283.8,
  283.9,     283.9,   283.9,   283.9,
  284.1,     284.1,   284.1,   284.1,
  284.45,    284.45,  284.45,  284.45,
  284.6,     284.6,   284.6,   284.6,
  284.65,    284.65,  284.65,  284.65,
  284.85,    284.85,  284.85,  284.85,
  284.9,     284.9,   284.9,   284.9,
  284.65,    284.65,  284.65,  284.65,
  284.5,     284.5,   284.5,   284.5,
  284.2,     284.2,   284.2,   284.2,
  283.55,    283.55,  283.55,  283.55,
  282.65,    282.65,  282.65,  282.65,
  281.95,    281.95,  281.95,  281.95,
  281.4,     281.4,   281.4,   281.4,
  280.7,     280.7,   280.7,   280.7,
  280.25,    280.25,  280.25,  280.25,
  279.75,    279.75,  279.75,  279.75,
  279.3,     279.3,   279.3,   279.3,
  279.35,    279.35,  279.35,  279.35,
  279.3,     279.3,   279.3,   279.3,
  278.65,    278.65,  278.65,  278.65,
  277.75,    277.75,  277.75,  277.75,
  277.4,     277.4,   277.4,   277.4,
  277.3,     277.3,   277.3,   277.3,
  277.05,    277.05,  277.05,  277.05,
  276.9,     276.9,   276.9,   276.9,
  277,       277,     277,     277,
  277.45,    277.45,  277.45,  277.45,
  277.9,     277.9,   277.9,   277.9,
  278.05,    278.05,  278.05,  278.05,
  277.95,    277.95,  277.95,  277.95,
  277.8,     277.8,   277.8,   277.8,
  278,       278,     278,     278,
  278.65,    278.65,  278.65,  278.65,
  279.35,    279.35,  279.35,  279.35,
  280.05,    280.05,  280.05,  280.05,
  280.9,     280.9,   280.9,   280.9,
  281.95,    281.95,  281.95,  281.95,
  283,       283,     283,     283,
  283.55,    283.55,  283.55,  283.55,
  283.85,    283.85,  283.85,  283.85,
  284.55,    284.55,  284.55,  284.55,
  285.5,     285.5,   285.5,   285.5,
  286.05,    286.05,  286.05,  286.05,
  286.35,    286.35,  286.35,  286.35,
  286.65,    286.65,  286.65,  286.65,
  286.8,     286.8,   286.8,   286.8,
  286.85,    286.85,  286.85,  286.85,
  286.85,    286.85,  286.85,  286.85,
  287,       287,     287,     287,
  287.25,    287.25,  287.25,  287.25,
  287.5,     287.5,   287.5,   287.5,
  287.75,    287.75,  287.75,  287.75,
  287.8,     287.8,   287.8,   287.8,
  287.75,    287.75,  287.75,  287.75,
  287.65,    287.65,  287.65,  287.65,
  287.35,    287.35,  287.35,  287.35,
  286.7,     286.7,   286.7,   286.7,
  285.95,    285.95,  285.95,  285.95,
  285.4,     285.4,   285.4,   285.4,
  284.95,    284.95,  284.95,  284.95,
  284.4,     284.4,   284.4,   284.4,
  283.9,     283.9,   283.9,   283.9,
  283.65,    283.65,  283.65,  283.65,
  283.25,    283.25,  283.25,  283.25,
  282.75,    282.75,  282.75,  282.75,
  282.5,     282.5,   282.5,   282.5,
  282.35,    282.35,  282.35,  282.35,
  282,       282,     282,     282,
  281.6,     281.6,   281.6,   281.6,
  281.5,     281.5,   281.5,   281.5,
  281.55,    281.55,  281.55,  281.55,
  281.45,    281.45,  281.45,  281.45,
  281.3,     281.3,   281.3,   281.3,
  281.1,     281.1,   281.1,   281.1,
  280.9,     280.9,   280.9,   280.9,
  280.75,    280.75,  280.75,  280.75,
  280.5,     280.5,   280.5,   280.5,
  280.25,    280.25,  280.25,  280.25,
  280.15,    280.15,  280.15,  280.15,
  280.25,    280.25,  280.25,  280.25,
  280.55,    280.55,  280.55,  280.55,
  281,       281,     281,     281,
  281.35,    281.35,  281.35,  281.35,
  281.65,    281.65,  281.65,  281.65,
  282.2,     282.2,   282.2,   282.2,
  282.8,     282.8,   282.8,   282.8,
  283.3,     283.3,   283.3,   283.3,
  283.75,    283.75,  283.75,  283.75,
  284.05,    284.05,  284.05,  284.05,
  284.2,     284.2,   284.2,   284.2,
  284.3,     284.3,   284.3,   284.3,
  284.4,     284.4,   284.4,   284.4,
  284.55,    284.55,  284.55,  284.55,
  284.2,     284.2,   284.2,   284.2,
  283.65,    283.65,  283.65,  283.65,
  283.55,    283.55,  283.55,  283.55,
  283.45,    283.45,  283.45,  283.45,
  283.1,     283.1,   283.1,   283.1,
  282.85,    282.85,  282.85,  282.85,
  282.95,    282.95,  282.95,  282.95,
  283.2,     283.2,   283.2,   283.2,
  283.35,    283.35,  283.35,  283.35,
  283.3,     283.3,   283.3,   283.3,
  283.2,     283.2,   283.2,   283.2,
  283,       283,     283,     283,
  282.75,    282.75,  282.75,  282.75,
  282.5,     282.5,   282.5,   282.5,
  282.2,     282.2,   282.2,   282.2,
  282,       282,     282,     282,
  281.85,    281.85,  281.85,  281.85,
  281.65,    281.65,  281.65,  281.65,
  281.45,    281.45,  281.45,  281.45,
  281.2,     281.2,   281.2,   281.2,
  280.95,    280.95,  280.95,  280.95,
  280.75,    280.75,  280.75,  280.75,
  280.65,    280.65,  280.65,  280.65,
  280.65,    280.65,  280.65,  280.65,
  280.6,     280.6,   280.6,   280.6,
  280.45,    280.45,  280.45,  280.45,
  280.25,    280.25,  280.25,  280.25,
  280.05,    280.05,  280.05,  280.05,
  280,       280,     280,     280,
  279.95,    279.95,  279.95,  279.95,
  279.65,    279.65,  279.65,  279.65,
  279.4,     279.4,   279.4,   279.4,
  279.35,    279.35,  279.35,  279.35,
  279.35,    279.35,  279.35,  279.35,
  279.4,     279.4,   279.4,   279.4,
  279.55,    279.55,  279.55,  279.55,
  279.85,    279.85,  279.85,  279.85,
  280.45,    280.45,  280.45,  280.45,
  281.2,     281.2,   281.2,   281.2,
  281.95,    281.95,  281.95,  281.95,
  282.65,    282.65,  282.65,  282.65,
  283.35,    283.35,  283.35,  283.35,
  284.1,     284.1,   284.1,   284.1,
  284.65,    284.65,  284.65,  284.65,
  284.95,    284.95,  284.95,  284.95,
  285.25,    285.25,  285.25,  285.25,
  285.7,     285.7,   285.7,   285.7,
  286,       286,     286,     286,
  286.35,    286.35,  286.35,  286.35,
  286.65,    286.65,  286.65,  286.65,
  286.85,    286.85,  286.85,  286.85,
  287.1,     287.1,   287.1,   287.1,
  287,       287,     287,     287,
  287,       287,     287,     287,
  287.3,     287.3,   287.3,   287.3,
  287.35,    287.35,  287.35,  287.35,
  287.2,     287.2,   287.2,   287.2,
  287.1,     287.1,   287.1,   287.1,
  286.95,    286.95,  286.95,  286.95,
  286.75,    286.75,  286.75,  286.75,
  286.55,    286.55,  286.55,  286.55,
  286.25,    286.25,  286.25,  286.25,
  285.95,    285.95,  285.95,  285.95,
  285.7,     285.7,   285.7,   285.7,
  284.95,    284.95,  284.95,  284.95,
  283.95,    283.95,  283.95,  283.95,
  283.45,    283.45,  283.45,  283.45,
  283.25,    283.25,  283.25,  283.25,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  283.1,     283.1,   283.1,   283.1,
  283.05,    283.05,  283.05,  283.05,
  282.95,    282.95,  282.95,  282.95,
  282.8,     282.8,   282.8,   282.8,
  282.7,     282.7,   282.7,   282.7,
  282.65,    282.65,  282.65,  282.65,
  282.6,     282.6,   282.6,   282.6,
  282.55,    282.55,  282.55,  282.55,
  282.6,     282.6,   282.6,   282.6,
  282.65,    282.65,  282.65,  282.65,
  282.65,    282.65,  282.65,  282.65,
  282.6,     282.6,   282.6,   282.6,
  282.55,    282.55,  282.55,  282.55,
  282.6,     282.6,   282.6,   282.6,
  282.65,    282.65,  282.65,  282.65,
  282.7,     282.7,   282.7,   282.7,
  282.85,    282.85,  282.85,  282.85,
  283,       283,     283,     283,
  283.2,     283.2,   283.2,   283.2,
  283.55,    283.55,  283.55,  283.55,
  283.95,    283.95,  283.95,  283.95,
  284.5,     284.5,   284.5,   284.5,
  285.05,    285.05,  285.05,  285.05,
  285.35,    285.35,  285.35,  285.35,
  285.75,    285.75,  285.75,  285.75,
  286.3,     286.3,   286.3,   286.3,
  286.55,    286.55,  286.55,  286.55,
  286.55,    286.55,  286.55,  286.55,
  286.8,     286.8,   286.8,   286.8,
  287.15,    287.15,  287.15,  287.15,
  286.8,     286.8,   286.8,   286.8,
  285.9,     285.9,   285.9,   285.9,
  285.35,    285.35,  285.35,  285.35,
  285.6,     285.6,   285.6,   285.6,
  286.25,    286.25,  286.25,  286.25,
  286.7,     286.7,   286.7,   286.7,
  286.9,     286.9,   286.9,   286.9,
  286.8,     286.8,   286.8,   286.8,
  286.3,     286.3,   286.3,   286.3,
  285.85,    285.85,  285.85,  285.85,
  285.55,    285.55,  285.55,  285.55,
  285,       285,     285,     285,
  284.45,    284.45,  284.45,  284.45,
  284.2,     284.2,   284.2,   284.2,
  284,       284,     284,     284,
  283.5,     283.5,   283.5,   283.5,
  282.9,     282.9,   282.9,   282.9,
  282.7,     282.7,   282.7,   282.7,
  282.8,     282.8,   282.8,   282.8,
  282.9,     282.9,   282.9,   282.9,
  283.05,    283.05,  283.05,  283.05,
  283.15,    283.15,  283.15,  283.15,
  283,       283,     283,     283,
  282.85,    282.85,  282.85,  282.85,
  282.85,    282.85,  282.85,  282.85,
  282.85,    282.85,  282.85,  282.85,
  282.75,    282.75,  282.75,  282.75,
  282.55,    282.55,  282.55,  282.55,
  282.2,     282.2,   282.2,   282.2,
  281.9,     281.9,   281.9,   281.9,
  281.95,    281.95,  281.95,  281.95,
  282.15,    282.15,  282.15,  282.15,
  282.55,    282.55,  282.55,  282.55,
  282.75,    282.75,  282.75,  282.75,
  282.55,    282.55,  282.55,  282.55,
  282.55,    282.55,  282.55,  282.55,
  282.8,     282.8,   282.8,   282.8,
  283.1,     283.1,   283.1,   283.1,
  283.4,     283.4,   283.4,   283.4,
  283.75,    283.75,  283.75,  283.75,
  284.1,     284.1,   284.1,   284.1,
  284.35,    284.35,  284.35,  284.35,
  284.55,    284.55,  284.55,  284.55,
  284.8,     284.8,   284.8,   284.8,
  285,       285,     285,     285,
  285.1,     285.1,   285.1,   285.1,
  285.45,    285.45,  285.45,  285.45,
  285.95,    285.95,  285.95,  285.95,
  286.15,    286.15,  286.15,  286.15,
  286.2,     286.2,   286.2,   286.2,
  286.45,    286.45,  286.45,  286.45,
  287,       287,     287,     287,
  287.35,    287.35,  287.35,  287.35,
  287.25,    287.25,  287.25,  287.25,
  287.05,    287.05,  287.05,  287.05,
  286.8,     286.8,   286.8,   286.8,
  285.95,    285.95,  285.95,  285.95,
  284.15,    284.15,  284.15,  284.15,
  282.9,     282.9,   282.9,   282.9,
  282.9,     282.9,   282.9,   282.9,
  283.25,    283.25,  283.25,  283.25,
  283.4,     283.4,   283.4,   283.4,
  283.35,    283.35,  283.35,  283.35,
  283.3,     283.3,   283.3,   283.3,
  283.3,     283.3,   283.3,   283.3,
  283.35,    283.35,  283.35,  283.35,
  283.35,    283.35,  283.35,  283.35,
  283.4,     283.4,   283.4,   283.4,
  283.45,    283.45,  283.45,  283.45,
  283.5,     283.5,   283.5,   283.5,
  283.55,    283.55,  283.55,  283.55,
  283.5,     283.5,   283.5,   283.5,
  283.4,     283.4,   283.4,   283.4,
  283.3,     283.3,   283.3,   283.3,
  283.1,     283.1,   283.1,   283.1,
  282.85,    282.85,  282.85,  282.85,
  282.7,     282.7,   282.7,   282.7,
  282.6,     282.6,   282.6,   282.6,
  282.55,    282.55,  282.55,  282.55,
  282.5,     282.5,   282.5,   282.5,
  282.5,     282.5,   282.5,   282.5,
  282.55,    282.55,  282.55,  282.55,
  282.45,    282.45,  282.45,  282.45,
  282.3,     282.3,   282.3,   282.3,
  282.15,    282.15,  282.15,  282.15,
  282,       282,     282,     282,
  281.95,    281.95,  281.95,  281.95,
  282,       282,     282,     282,
  282.1,     282.1,   282.1,   282.1,
  282.2,     282.2,   282.2,   282.2,
  282.25,    282.25,  282.25,  282.25,
  282.15,    282.15,  282.15,  282.15,
  282.05,    282.05,  282.05,  282.05,
  282.1,     282.1,   282.1,   282.1,
  282.2,     282.2,   282.2,   282.2,
  282.4,     282.4,   282.4,   282.4,
  282.7,     282.7,   282.7,   282.7,
  282.9,     282.9,   282.9,   282.9,
  282.95,    282.95,  282.95,  282.95,
  282.95,    282.95,  282.95,  282.95,
  282.9,     282.9,   282.9,   282.9,
  282.75,    282.75,  282.75,  282.75,
  282.55,    282.55,  282.55,  282.55,
  282.5,     282.5,   282.5,   282.5,
  282.5,     282.5,   282.5,   282.5,
  282.15,    282.15,  282.15,  282.15,
  281.65,    281.65,  281.65,  281.65,
  281.4,     281.4,   281.4,   281.4,
  281.3,     281.3,   281.3,   281.3,
  281.25,    281.25,  281.25,  281.25,
  281.25,    281.25,  281.25,  281.25,
  281.25,    281.25,  281.25,  281.25,
  281.3,     281.3,   281.3,   281.3,
  281.35,    281.35,  281.35,  281.35,
  281.35,    281.35,  281.35,  281.35,
  281.4,     281.4,   281.4,   281.4,
  281.3,     281.3,   281.3,   281.3,
  281,       281,     281,     281,
  280.7,     280.7,   280.7,   280.7,
  280.4,     280.4,   280.4,   280.4,
  280.2,     280.2,   280.2,   280.2,
  280.05,    280.05,  280.05,  280.05,
  279.8,     279.8,   279.8,   279.8,
  279.65,    279.65,  279.65,  279.65,
  279.55,    279.55,  279.55,  279.55,
  279.45,    279.45,  279.45,  279.45,
  279.75,    279.75,  279.75,  279.75,
  280.25,    280.25,  280.25,  280.25,
  280.5,     280.5,   280.5,   280.5,
  280.85,    280.85,  280.85,  280.85,
  281.4,     281.4,   281.4,   281.4,
  281.75,    281.75,  281.75,  281.75,
  281.95,    281.95,  281.95,  281.95,
  282.05,    282.05,  282.05,  282.05,
  282.2,     282.2,   282.2,   282.2,
  282.85,    282.85,  282.85,  282.85,
  283.85,    283.85,  283.85,  283.85,
  284.7,     284.7,   284.7,   284.7,
  285.2,     285.2,   285.2,   285.2,
  285.25,    285.25,  285.25,  285.25,
  285.25,    285.25,  285.25,  285.25,
  285.55,    285.55,  285.55,  285.55,
  285.75,    285.75,  285.75,  285.75,
  285.8,     285.8,   285.8,   285.8,
  285.75,    285.75,  285.75,  285.75,
  285.6,     285.6,   285.6,   285.6,
  285.4,     285.4,   285.4,   285.4,
  285,       285,     285,     285,
  284.5,     284.5,   284.5,   284.5,
  284.2,     284.2,   284.2,   284.2,
  284.1,     284.1,   284.1,   284.1,
  284.15,    284.15,  284.15,  284.15,
  284.2,     284.2,   284.2,   284.2,
  284.1,     284.1,   284.1,   284.1,
  283.85,    283.85,  283.85,  283.85,
  283.5,     283.5,   283.5,   283.5,
  283.15,    283.15,  283.15,  283.15,
  282.7,     282.7,   282.7,   282.7,
  282.15,    282.15,  282.15,  282.15,
  281.8,     281.8,   281.8,   281.8,
  281.55,    281.55,  281.55,  281.55,
  281.15,    281.15,  281.15,  281.15,
  280.6,     280.6,   280.6,   280.6,
  280.2,     280.2,   280.2,   280.2,
  279.8,     279.8,   279.8,   279.8,
  279.3,     279.3,   279.3,   279.3,
  279.1,     279.1,   279.1,   279.1,
  278.8,     278.8,   278.8,   278.8,
  278.2,     278.2,   278.2,   278.2,
  277.55,    277.55,  277.55,  277.55,
  277.05,    277.05,  277.05,  277.05,
  276.55,    276.55,  276.55,  276.55,
  276.05,    276.05,  276.05,  276.05,
  275.95,    275.95,  275.95,  275.95,
  276.15,    276.15,  276.15,  276.15,
  277,       277,     277,     277,
  278.6,     278.6,   278.6,   278.6,
  280.15,    280.15,  280.15,  280.15,
  281.3,     281.3,   281.3,   281.3,
  282.15,    282.15,  282.15,  282.15,
  283.2,     283.2,   283.2,   283.2,
  284.5,     284.5,   284.5,   284.5,
  285.6,     285.6,   285.6,   285.6,
  286.5,     286.5,   286.5,   286.5,
  287.1,     287.1,   287.1,   287.1,
  287.45,    287.45,  287.45,  287.45,
  287.8,     287.8,   287.8,   287.8,
  288.35,    288.35,  288.35,  288.35,
  288.85,    288.85,  288.85,  288.85,
  289.3,     289.3,   289.3,   289.3,
  290.1,     290.1,   290.1,   290.1,
  290.6,     290.6,   290.6,   290.6,
  290.5,     290.5,   290.5,   290.5,
  290.45,    290.45,  290.45,  290.45,
  290.55,    290.55,  290.55,  290.55,
  290.65,    290.65,  290.65,  290.65,
  290.8,     290.8,   290.8,   290.8,
  290.9,     290.9,   290.9,   290.9,
  291,       291,     291,     291,
  290.9,     290.9,   290.9,   290.9,
  290.45,    290.45,  290.45,  290.45,
  289.75,    289.75,  289.75,  289.75,
  288.75,    288.75,  288.75,  288.75,
  287.65,    287.65,  287.65,  287.65,
  286.8,     286.8,   286.8,   286.8,
  286.1,     286.1,   286.1,   286.1,
  285.35,    285.35,  285.35,  285.35,
  284.8,     284.8,   284.8,   284.8,
  284.55,    284.55,  284.55,  284.55,
  284.4,     284.4,   284.4,   284.4,
  284.4,     284.4,   284.4,   284.4,
  284.35,    284.35,  284.35,  284.35,
  284,       284,     284,     284,
  283.65,    283.65,  283.65,  283.65,
  283.5,     283.5,   283.5,   283.5,
  283.4,     283.4,   283.4,   283.4,
  283.1,     283.1,   283.1,   283.1,
  282.45,    282.45,  282.45,  282.45,
  281.8,     281.8,   281.8,   281.8,
  281.2,     281.2,   281.2,   281.2,
  280.8,     280.8,   280.8,   280.8,
  280.7,     280.7,   280.7,   280.7,
  280.8,     280.8,   280.8,   280.8,
  281.4,     281.4,   281.4,   281.4,
  282.7,     282.7,   282.7,   282.7,
  284.5,     284.5,   284.5,   284.5,
  286.1,     286.1,   286.1,   286.1,
  287.5,     287.5,   287.5,   287.5,
  288.75,    288.75,  288.75,  288.75,
  289.5,     289.5,   289.5,   289.5,
  290.05,    290.05,  290.05,  290.05,
  290.75,    290.75,  290.75,  290.75,
  291.4,     291.4,   291.4,   291.4,
  291.9,     291.9,   291.9,   291.9,
  292.45,    292.45,  292.45,  292.45,
  293.1,     293.1,   293.1,   293.1,
  293.6,     293.6,   293.6,   293.6,
  294.05,    294.05,  294.05,  294.05,
  294.4,     294.4,   294.4,   294.4,
  294.5,     294.5,   294.5,   294.5,
  294.6,     294.6,   294.6,   294.6,
  294.75,    294.75,  294.75,  294.75,
  294.9,     294.9,   294.9,   294.9,
  295.15,    295.15,  295.15,  295.15,
  295.2,     295.2,   295.2,   295.2,
  294.9,     294.9,   294.9,   294.9,
  294.55,    294.55,  294.55,  294.55,
  293.95,    293.95,  293.95,  293.95,
  293,       293,     293,     293,
  291.8,     291.8,   291.8,   291.8,
  290.5,     290.5,   290.5,   290.5,
  289.45,    289.45,  289.45,  289.45,
  288.8,     288.8,   288.8,   288.8,
  288.3,     288.3,   288.3,   288.3,
  288,       288,     288,     288,
  287.35,    287.35,  287.35,  287.35,
  286.9,     286.9,   286.9,   286.9,
  286.65,    286.65,  286.65,  286.65,
  285.55,    285.55,  285.55,  285.55,
  284.65,    284.65,  284.65,  284.65,
  283.85,    283.85,  283.85,  283.85,
  282.7,     282.7,   282.7,   282.7,
  283,       283,     283,     283,
  283.6,     283.6,   283.6,   283.6,
  283.2,     283.2,   283.2,   283.2,
  282.8,     282.8,   282.8,   282.8,
  282.55,    282.55,  282.55,  282.55,
  282.45,    282.45,  282.45,  282.45,
  282.1,     282.1,   282.1,   282.1,
  282.2,     282.2,   282.2,   282.2,
  282.7,     282.7,   282.7,   282.7,
  283.2,     283.2,   283.2,   283.2,
  284.05,    284.05,  284.05,  284.05,
  285.15,    285.15,  285.15,  285.15,
  286.45,    286.45,  286.45,  286.45,
  287.6,     287.6,   287.6,   287.6,
  288.4,     288.4,   288.4,   288.4,
  289.2,     289.2,   289.2,   289.2,
  290,       290,     290,     290,
  290.6,     290.6,   290.6,   290.6,
  291.15,    291.15,  291.15,  291.15,
  291.6,     291.6,   291.6,   291.6,
  292,       292,     292,     292,
  292.5,     292.5,   292.5,   292.5,
  293.05,    293.05,  293.05,  293.05,
  293.65,    293.65,  293.65,  293.65,
  294.05,    294.05,  294.05,  294.05,
  294.45,    294.45,  294.45,  294.45,
  294.9,     294.9,   294.9,   294.9,
  295.15,    295.15,  295.15,  295.15,
  295,       295,     295,     295,
  294.65,    294.65,  294.65,  294.65,
  294.25,    294.25,  294.25,  294.25,
  293.65,    293.65,  293.65,  293.65,
  292.9,     292.9,   292.9,   292.9,
  292.1,     292.1,   292.1,   292.1,
  291.4,     291.4,   291.4,   291.4,
  290.65,    290.65,  290.65,  290.65,
  290,       290,     290,     290,
  289.55,    289.55,  289.55,  289.55,
  289.2,     289.2,   289.2,   289.2,
  288.95,    288.95,  288.95,  288.95,
  288.7,     288.7,   288.7,   288.7,
  288.45,    288.45,  288.45,  288.45,
  288.25,    288.25,  288.25,  288.25,
  288,       288,     288,     288,
  287.75,    287.75,  287.75,  287.75,
  287.55,    287.55,  287.55,  287.55,
  287.3,     287.3,   287.3,   287.3,
  287,       287,     287,     287,
  286.8,     286.8,   286.8,   286.8,
  286.6,     286.6,   286.6,   286.6,
  286.3,     286.3,   286.3,   286.3,
  286.15,    286.15,  286.15,  286.15,
  286.2,     286.2,   286.2,   286.2,
  286.45,    286.45,  286.45,  286.45,
  286.6,     286.6,   286.6,   286.6,
  286.45,    286.45,  286.45,  286.45,
  286.4,     286.4,   286.4,   286.4,
  286.35,    286.35,  286.35,  286.35,
  286.25,    286.25,  286.25,  286.25,
  286.25,    286.25,  286.25,  286.25,
  286.1,     286.1,   286.1,   286.1,
  285.95,    285.95,  285.95,  285.95,
  285.95,    285.95,  285.95,  285.95,
  286.25,    286.25,  286.25,  286.25,
  287.15,    287.15,  287.15,  287.15,
  288.25,    288.25,  288.25,  288.25,
  288.65,    288.65,  288.65,  288.65,
  288.95,    288.95,  288.95,  288.95,
  289.8,     289.8,   289.8,   289.8,
  290.45,    290.45,  290.45,  290.45,
  290.6,     290.6,   290.6,   290.6,
  290.7,     290.7,   290.7,   290.7,
  290.9,     290.9,   290.9,   290.9,
  290.5,     290.5,   290.5,   290.5,
  289.45,    289.45,  289.45,  289.45,
  289.15,    289.15,  289.15,  289.15,
  288.9,     288.9,   288.9,   288.9,
  288.2,     288.2,   288.2,   288.2,
  288,       288,     288,     288,
  287.9,     287.9,   287.9,   287.9,
  287.8,     287.8,   287.8,   287.8,
  287.85,    287.85,  287.85,  287.85,
  288,       288,     288,     288,
  288.05,    288.05,  288.05,  288.05,
  288.15,    288.15,  288.15,  288.15,
  288.3,     288.3,   288.3,   288.3,
  288.4,     288.4,   288.4,   288.4,
  288.25,    288.25,  288.25,  288.25,
  287.75,    287.75,  287.75,  287.75,
  287.15,    287.15,  287.15,  287.15,
  286.6,     286.6,   286.6,   286.6,
  286.15,    286.15,  286.15,  286.15,
  285.9,     285.9,   285.9,   285.9,
  285.8,     285.8,   285.8,   285.8,
  285.6,     285.6,   285.6,   285.6,
  285.15,    285.15,  285.15,  285.15,
  284.7,     284.7,   284.7,   284.7,
  284.65,    284.65,  284.65,  284.65,
  284.85,    284.85,  284.85,  284.85,
  285.1,     285.1,   285.1,   285.1,
  285.2,     285.2,   285.2,   285.2,
  285.15,    285.15,  285.15,  285.15,
  285.15,    285.15,  285.15,  285.15,
  285.2,     285.2,   285.2,   285.2,
  285.35,    285.35,  285.35,  285.35,
  285.6,     285.6,   285.6,   285.6,
  285.8,     285.8,   285.8,   285.8,
  285.9,     285.9,   285.9,   285.9,
  286.05,    286.05,  286.05,  286.05,
  285.6,     285.6,   285.6,   285.6,
  285.05,    285.05,  285.05,  285.05,
  285.75,    285.75,  285.75,  285.75,
  286.65,    286.65,  286.65,  286.65,
  287,       287,     287,     287,
  287.25,    287.25,  287.25,  287.25,
  287.6,     287.6,   287.6,   287.6,
  287.8,     287.8,   287.8,   287.8,
  288.15,    288.15,  288.15,  288.15,
  288.65,    288.65,  288.65,  288.65,
  287.6,     287.6,   287.6,   287.6,
  285.5,     285.5,   285.5,   285.5,
  284.35,    284.35,  284.35,  284.35,
  284.4,     284.4,   284.4,   284.4,
  284.85,    284.85,  284.85,  284.85,
  285.45,    285.45,  285.45,  285.45,
  286.05,    286.05,  286.05,  286.05,
  286.4,     286.4,   286.4,   286.4,
  286.65,    286.65,  286.65,  286.65,
  286.75,    286.75,  286.75,  286.75,
  286.75,    286.75,  286.75,  286.75,
  286.65,    286.65,  286.65,  286.65,
  286.4,     286.4,   286.4,   286.4,
  286,       286,     286,     286,
  285.45,    285.45,  285.45,  285.45,
  285,       285,     285,     285,
  284.8,     284.8,   284.8,   284.8,
  284.85,    284.85,  284.85,  284.85,
  285,       285,     285,     285,
  285.05,    285.05,  285.05,  285.05,
  284.95,    284.95,  284.95,  284.95,
  284.75,    284.75,  284.75,  284.75,
  284.55,    284.55,  284.55,  284.55,
  284.45,    284.45,  284.45,  284.45,
  284.65,    284.65,  284.65,  284.65,
  284.95,    284.95,  284.95,  284.95,
  284.8,     284.8,   284.8,   284.8,
  284.15,    284.15,  284.15,  284.15,
  283.7,     283.7,   283.7,   283.7,
  283.8,     283.8,   283.8,   283.8,
  284.05,    284.05,  284.05,  284.05,
  284.2,     284.2,   284.2,   284.2,
  284.2,     284.2,   284.2,   284.2,
  283.35,    283.35,  283.35,  283.35,
  281.7,     281.7,   281.7,   281.7,
  280.35,    280.35,  280.35,  280.35,
  279.6,     279.6,   279.6,   279.6,
  279.15,    279.15,  279.15,  279.15,
  278.85,    278.85,  278.85,  278.85,
  278.65,    278.65,  278.65,  278.65,
  278.55,    278.55,  278.55,  278.55,
  278.6,     278.6,   278.6,   278.6,
  278.6,     278.6,   278.6,   278.6,
  278.65,    278.65,  278.65,  278.65,
  278.65,    278.65,  278.65,  278.65,
  278.45,    278.45,  278.45,  278.45,
  278.2,     278.2,   278.2,   278.2,
  277.85,    277.85,  277.85,  277.85,
  277.6,     277.6,   277.6,   277.6,
  277.6,     277.6,   277.6,   277.6,
  277.65,    277.65,  277.65,  277.65,
  277.8,     277.8,   277.8,   277.8,
  277.9,     277.9,   277.9,   277.9,
  278,       278,     278,     278,
  278.25,    278.25,  278.25,  278.25,
  278.65,    278.65,  278.65,  278.65,
  278.9,     278.9,   278.9,   278.9,
  279.05,    279.05,  279.05,  279.05,
  279.2,     279.2,   279.2,   279.2,
  279.05,    279.05,  279.05,  279.05,
  278.7,     278.7,   278.7,   278.7,
  278,       278,     278,     278,
  277.05,    277.05,  277.05,  277.05,
  276.55,    276.55,  276.55,  276.55,
  276.5,     276.5,   276.5,   276.5,
  276.35,    276.35,  276.35,  276.35,
  276.05,    276.05,  276.05,  276.05,
  275.8,     275.8,   275.8,   275.8,
  275.7,     275.7,   275.7,   275.7,
  275.6,     275.6,   275.6,   275.6,
  275.4,     275.4,   275.4,   275.4,
  275.2,     275.2,   275.2,   275.2,
  274.8,     274.8,   274.8,   274.8,
  274.4,     274.4,   274.4,   274.4,
  274.35,    274.35,  274.35,  274.35,
  274.45,    274.45,  274.45,  274.45,
  274.2,     274.2,   274.2,   274.2,
  273.75,    273.75,  273.75,  273.75,
  273.5,     273.5,   273.5,   273.5,
  273.25,    273.25,  273.25,  273.25,
  273.3,     273.3,   273.3,   273.3,
  274.05,    274.05,  274.05,  274.05,
  275.25,    275.25,  275.25,  275.25,
  276.35,    276.35,  276.35,  276.35,
  277.4,     277.4,   277.4,   277.4,
  278.45,    278.45,  278.45,  278.45,
  279.25,    279.25,  279.25,  279.25,
  279.6,     279.6,   279.6,   279.6,
  279.8,     279.8,   279.8,   279.8,
  280.1,     280.1,   280.1,   280.1,
  279.1,     279.1,   279.1,   279.1,
  278.45,    278.45,  278.45,  278.45,
  279.35,    279.35,  279.35,  279.35,
  280.2,     280.2,   280.2,   280.2,
  280.5,     280.5,   280.5,   280.5,
  279.5,     279.5,   279.5,   279.5,
  278.65,    278.65,  278.65,  278.65,
  278.5,     278.5,   278.5,   278.5,
  278.75,    278.75,  278.75,  278.75,
  279.35,    279.35,  279.35,  279.35,
  279.95,    279.95,  279.95,  279.95,
  280.85,    280.85,  280.85,  280.85,
  281.1,     281.1,   281.1,   281.1,
  281,       281,     281,     281,
  281.25,    281.25,  281.25,  281.25,
  281.45,    281.45,  281.45,  281.45,
  281.65,    281.65,  281.65,  281.65,
  281.7,     281.7,   281.7,   281.7,
  281.4,     281.4,   281.4,   281.4,
  280.75,    280.75,  280.75,  280.75,
  279.8,     279.8,   279.8,   279.8,
  278.9,     278.9,   278.9,   278.9,
  278.35,    278.35,  278.35,  278.35,
  278.1,     278.1,   278.1,   278.1,
  277.9,     277.9,   277.9,   277.9,
  277.55,    277.55,  277.55,  277.55,
  277.2,     277.2,   277.2,   277.2,
  276.8,     276.8,   276.8,   276.8,
  276.35,    276.35,  276.35,  276.35,
  276.05,    276.05,  276.05,  276.05,
  275.8,     275.8,   275.8,   275.8,
  275.6,     275.6,   275.6,   275.6,
  275.55,    275.55,  275.55,  275.55,
  275.4,     275.4,   275.4,   275.4,
  275.1,     275.1,   275.1,   275.1,
  274.9,     274.9,   274.9,   274.9,
  274.8,     274.8,   274.8,   274.8,
  274.75,    274.75,  274.75,  274.75,
  274.95,    274.95,  274.95,  274.95,
  275.55,    275.55,  275.55,  275.55,
  276.45,    276.45,  276.45,  276.45,
  277.5,     277.5,   277.5,   277.5,
  278.65,    278.65,  278.65,  278.65,
  279.7,     279.7,   279.7,   279.7,
  280.35,    280.35,  280.35,  280.35,
  280.6,     280.6,   280.6,   280.6,
  280.9,     280.9,   280.9,   280.9,
  281.35,    281.35,  281.35,  281.35,
  281.8,     281.8,   281.8,   281.8,
  281.85,    281.85,  281.85,  281.85,
  281.3,     281.3,   281.3,   281.3,
  281,       281,     281,     281,
  280.55,    280.55,  280.55,  280.55,
  280,       280,     280,     280,
  280.3,     280.3,   280.3,   280.3,
  280.95,    280.95,  280.95,  280.95,
  281.45,    281.45,  281.45,  281.45,
  281.9,     281.9,   281.9,   281.9,
  282.35,    282.35,  282.35,  282.35,
  282.8,     282.8,   282.8,   282.8,
  282.5,     282.5,   282.5,   282.5,
  281.2,     281.2,   281.2,   281.2,
  280.45,    280.45,  280.45,  280.45,
  280.65,    280.65,  280.65,  280.65,
  280.95,    280.95,  280.95,  280.95,
  281.1,     281.1,   281.1,   281.1,
  281,       281,     281,     281,
  280.7,     280.7,   280.7,   280.7,
  280.55,    280.55,  280.55,  280.55,
  280.4,     280.4,   280.4,   280.4,
  280.15,    280.15,  280.15,  280.15,
  280.15,    280.15,  280.15,  280.15,
  280.3,     280.3,   280.3,   280.3,
  280.4,     280.4,   280.4,   280.4,
  280.6,     280.6,   280.6,   280.6,
  280.85,    280.85,  280.85,  280.85,
  280.8,     280.8,   280.8,   280.8,
  280.65,    280.65,  280.65,  280.65,
  280.55,    280.55,  280.55,  280.55,
  280.35,    280.35,  280.35,  280.35,
  280.3,     280.3,   280.3,   280.3,
  280.25,    280.25,  280.25,  280.25,
  279.8,     279.8,   279.8,   279.8,
  279.4,     279.4,   279.4,   279.4,
  279.35,    279.35,  279.35,  279.35,
  279.4,     279.4,   279.4,   279.4,
  279.6,     279.6,   279.6,   279.6,
  279.85,    279.85,  279.85,  279.85,
  280.1,     280.1,   280.1,   280.1,
  280.35,    280.35,  280.35,  280.35,
  280.75,    280.75,  280.75,  280.75,
  281.45,    281.45,  281.45,  281.45,
  281.9,     281.9,   281.9,   281.9,
  281.25,    281.25,  281.25,  281.25,
  281.05,    281.05,  281.05,  281.05,
  282.05,    282.05,  282.05,  282.05,
  282.35,    282.35,  282.35,  282.35,
  282.15,    282.15,  282.15,  282.15,
  282.3,     282.3,   282.3,   282.3,
  282.15,    282.15,  282.15,  282.15,
  282.45,    282.45,  282.45,  282.45,
  283.25,    283.25,  283.25,  283.25,
  283.45,    283.45,  283.45,  283.45,
  283.8,     283.8,   283.8,   283.8,
  283.7,     283.7,   283.7,   283.7,
  282.95,    282.95,  282.95,  282.95,
  282.45,    282.45,  282.45,  282.45,
  282.25,    282.25,  282.25,  282.25,
  282.3,     282.3,   282.3,   282.3,
  282.5,     282.5,   282.5,   282.5,
  282.85,    282.85,  282.85,  282.85,
  283.35,    283.35,  283.35,  283.35,
  283.7,     283.7,   283.7,   283.7,
  283.65,    283.65,  283.65,  283.65,
  283.15,    283.15,  283.15,  283.15,
  282.25,    282.25,  282.25,  282.25,
  281.5,     281.5,   281.5,   281.5,
  281.05,    281.05,  281.05,  281.05,
  280.7,     280.7,   280.7,   280.7,
  280.7,     280.7,   280.7,   280.7,
  281.1,     281.1,   281.1,   281.1,
  281.4,     281.4,   281.4,   281.4,
  281.3,     281.3,   281.3,   281.3,
  281.1,     281.1,   281.1,   281.1,
  281.05,    281.05,  281.05,  281.05,
  281.05,    281.05,  281.05,  281.05,
  281.1,     281.1,   281.1,   281.1,
  280.95,    280.95,  280.95,  280.95,
  280.55,    280.55,  280.55,  280.55,
  280.25,    280.25,  280.25,  280.25,
  280.2,     280.2,   280.2,   280.2,
  280.25,    280.25,  280.25,  280.25,
  280.25,    280.25,  280.25,  280.25,
  280.4,     280.4,   280.4,   280.4,
  280.75,    280.75,  280.75,  280.75,
  281,       281,     281,     281,
  281.1,     281.1,   281.1,   281.1,
  281.3,     281.3,   281.3,   281.3,
  281.6,     281.6,   281.6,   281.6,
  282.05,    282.05,  282.05,  282.05,
  282.8,     282.8,   282.8,   282.8,
  283.5,     283.5,   283.5,   283.5,
  284,       284,     284,     284,
  284.65,    284.65,  284.65,  284.65,
  285.35,    285.35,  285.35,  285.35,
  285.95,    285.95,  285.95,  285.95,
  285.25,    285.25,  285.25,  285.25,
  285.1,     285.1,   285.1,   285.1,
  286.1,     286.1,   286.1,   286.1,
  286.5,     286.5,   286.5,   286.5,
  287.15,    287.15,  287.15,  287.15,
  287.6,     287.6,   287.6,   287.6,
  287.5,     287.5,   287.5,   287.5,
  287.65,    287.65,  287.65,  287.65,
  287.95,    287.95,  287.95,  287.95,
  288,       288,     288,     288,
  288.25,    288.25,  288.25,  288.25,
  288.45,    288.45,  288.45,  288.45,
  288.3,     288.3,   288.3,   288.3,
  288.15,    288.15,  288.15,  288.15,
  288.2,     288.2,   288.2,   288.2,
  288.2,     288.2,   288.2,   288.2,
  287.95,    287.95,  287.95,  287.95,
  287.65,    287.65,  287.65,  287.65,
  287.45,    287.45,  287.45,  287.45,
  287.3,     287.3,   287.3,   287.3,
  286.7,     286.7,   286.7,   286.7,
  285.7,     285.7,   285.7,   285.7,
  285.25,    285.25,  285.25,  285.25,
  285.45,    285.45,  285.45,  285.45,
  285.55,    285.55,  285.55,  285.55,
  285.05,    285.05,  285.05,  285.05,
  284.55,    284.55,  284.55,  284.55,
  284.3,     284.3,   284.3,   284.3,
  284.15,    284.15,  284.15,  284.15,
  284.1,     284.1,   284.1,   284.1,
  284,       284,     284,     284,
  283.9,     283.9,   283.9,   283.9,
  283.8,     283.8,   283.8,   283.8,
  283.7,     283.7,   283.7,   283.7,
  283.65,    283.65,  283.65,  283.65,
  283.7,     283.7,   283.7,   283.7,
  283.75,    283.75,  283.75,  283.75,
  283.85,    283.85,  283.85,  283.85,
  284.15,    284.15,  284.15,  284.15,
  284.7,     284.7,   284.7,   284.7,
  285.15,    285.15,  285.15,  285.15,
  285.65,    285.65,  285.65,  285.65,
  286.3,     286.3,   286.3,   286.3,
  286.65,    286.65,  286.65,  286.65,
  286.9,     286.9,   286.9,   286.9,
  287,       287,     287,     287,
  287.2,     287.2,   287.2,   287.2,
  287.55,    287.55,  287.55,  287.55,
  287.85,    287.85,  287.85,  287.85,
  287.9,     287.9,   287.9,   287.9,
  287.95,    287.95,  287.95,  287.95,
  288.3,     288.3,   288.3,   288.3,
  288.45,    288.45,  288.45,  288.45,
  288.4,     288.4,   288.4,   288.4,
  288.45,    288.45,  288.45,  288.45,
  288.45,    288.45,  288.45,  288.45,
  287.75,    287.75,  287.75,  287.75,
  287.4,     287.4,   287.4,   287.4,
  288.3,     288.3,   288.3,   288.3,
  288.9,     288.9,   288.9,   288.9,
  288.2,     288.2,   288.2,   288.2,
  286.3,     286.3,   286.3,   286.3,
  284.4,     284.4,   284.4,   284.4,
  283.75,    283.75,  283.75,  283.75,
  283.8,     283.8,   283.8,   283.8,
  283.9,     283.9,   283.9,   283.9,
  284.05,    284.05,  284.05,  284.05,
  284.4,     284.4,   284.4,   284.4,
  284.7,     284.7,   284.7,   284.7,
  284.8,     284.8,   284.8,   284.8,
  284.9,     284.9,   284.9,   284.9,
  284.9,     284.9,   284.9,   284.9,
  284.85,    284.85,  284.85,  284.85,
  284.65,    284.65,  284.65,  284.65,
  284.45,    284.45,  284.45,  284.45,
  284.4,     284.4,   284.4,   284.4,
  284.2,     284.2,   284.2,   284.2,
  283.9,     283.9,   283.9,   283.9,
  283.5,     283.5,   283.5,   283.5,
  283,       283,     283,     283,
  282.75,    282.75,  282.75,  282.75,
  282.7,     282.7,   282.7,   282.7,
  282.6,     282.6,   282.6,   282.6,
  282.6,     282.6,   282.6,   282.6,
  282.75,    282.75,  282.75,  282.75,
  283.05,    283.05,  283.05,  283.05,
  283.45,    283.45,  283.45,  283.45,
  283.9,     283.9,   283.9,   283.9,
  284.4,     284.4,   284.4,   284.4,
  284.9,     284.9,   284.9,   284.9,
  285.15,    285.15,  285.15,  285.15,
  285.1,     285.1,   285.1,   285.1,
  284.95,    284.95,  284.95,  284.95,
  285.05,    285.05,  285.05,  285.05,
  285.45,    285.45,  285.45,  285.45,
  285.9,     285.9,   285.9,   285.9,
  286.4,     286.4,   286.4,   286.4,
  287.05,    287.05,  287.05,  287.05,
  287.35,    287.35,  287.35,  287.35,
  287.75,    287.75,  287.75,  287.75,
  288.45,    288.45,  288.45,  288.45,
  288.45,    288.45,  288.45,  288.45,
  288.55,    288.55,  288.55,  288.55,
  289,       289,     289,     289,
  289.2,     289.2,   289.2,   289.2,
  289.2,     289.2,   289.2,   289.2,
  289.45,    289.45,  289.45,  289.45,
  289.85,    289.85,  289.85,  289.85,
  289.75,    289.75,  289.75,  289.75,
  288.8,     288.8,   288.8,   288.8,
  287,       287,     287,     287,
  285.7,     285.7,   285.7,   285.7,
  285.4,     285.4,   285.4,   285.4,
  285.15,    285.15,  285.15,  285.15,
  284.7,     284.7,   284.7,   284.7,
  284.2,     284.2,   284.2,   284.2,
  283.9,     283.9,   283.9,   283.9,
  283.25,    283.25,  283.25,  283.25,
  282.35,    282.35,  282.35,  282.35,
  281.8,     281.8,   281.8,   281.8,
  281.55,    281.55,  281.55,  281.55,
  281.3,     281.3,   281.3,   281.3,
  280.95,    280.95,  280.95,  280.95,
  280.95,    280.95,  280.95,  280.95,
  281,       281,     281,     281,
  280.75,    280.75,  280.75,  280.75,
  280.4,     280.4,   280.4,   280.4,
  280.25,    280.25,  280.25,  280.25,
  280.2,     280.2,   280.2,   280.2,
  280.25,    280.25,  280.25,  280.25,
  280.4,     280.4,   280.4,   280.4,
  280.35,    280.35,  280.35,  280.35,
  280.5,     280.5,   280.5,   280.5,
  281.2,     281.2,   281.2,   281.2,
  282.2,     282.2,   282.2,   282.2,
  283.6,     283.6,   283.6,   283.6,
  285.3,     285.3,   285.3,   285.3,
  286.6,     286.6,   286.6,   286.6,
  287.3,     287.3,   287.3,   287.3,
  288,       288,     288,     288,
  288.8,     288.8,   288.8,   288.8,
  289.5,     289.5,   289.5,   289.5,
  290.15,    290.15,  290.15,  290.15,
  290.55,    290.55,  290.55,  290.55,
  290.55,    290.55,  290.55,  290.55,
  290.85,    290.85,  290.85,  290.85,
  291.35,    291.35,  291.35,  291.35,
  291.95,    291.95,  291.95,  291.95,
  292.3,     292.3,   292.3,   292.3,
  292.55,    292.55,  292.55,  292.55,
  292.85,    292.85,  292.85,  292.85,
  292.95,    292.95,  292.95,  292.95,
  293.2,     293.2,   293.2,   293.2,
  293.1,     293.1,   293.1,   293.1,
  292.8,     292.8,   292.8,   292.8,
  292.8,     292.8,   292.8,   292.8,
  292.65,    292.65,  292.65,  292.65,
  292.35,    292.35,  292.35,  292.35,
  292.2,     292.2,   292.2,   292.2,
  291.75,    291.75,  291.75,  291.75,
  291.2,     291.2,   291.2,   291.2,
  290.75,    290.75,  290.75,  290.75,
  290.15,    290.15,  290.15,  290.15,
  289.05,    289.05,  289.05,  289.05,
  288.15,    288.15,  288.15,  288.15,
  287.65,    287.65,  287.65,  287.65,
  287.05,    287.05,  287.05,  287.05,
  286.65,    286.65,  286.65,  286.65,
  286.4,     286.4,   286.4,   286.4,
  286.05,    286.05,  286.05,  286.05,
  285.8,     285.8,   285.8,   285.8,
  285.7,     285.7,   285.7,   285.7,
  285.7,     285.7,   285.7,   285.7,
  285.55,    285.55,  285.55,  285.55,
  285.4,     285.4,   285.4,   285.4,
  285.25,    285.25,  285.25,  285.25,
  284.6,     284.6,   284.6,   284.6,
  283.9,     283.9,   283.9,   283.9,
  283.95,    283.95,  283.95,  283.95,
  284.1,     284.1,   284.1,   284.1,
  283.9,     283.9,   283.9,   283.9,
  283.9,     283.9,   283.9,   283.9,
  284.1,     284.1,   284.1,   284.1,
  284.45,    284.45,  284.45,  284.45,
  284.75,    284.75,  284.75,  284.75,
  284.85,    284.85,  284.85,  284.85,
  284.9,     284.9,   284.9,   284.9,
  284.95,    284.95,  284.95,  284.95,
  284.9,     284.9,   284.9,   284.9,
  284.8,     284.8,   284.8,   284.8,
  284.75,    284.75,  284.75,  284.75,
  284.6,     284.6,   284.6,   284.6,
  284.4,     284.4,   284.4,   284.4,
  284.35,    284.35,  284.35,  284.35,
  284,       284,     284,     284,
  283.6,     283.6,   283.6,   283.6,
  283.5,     283.5,   283.5,   283.5,
  283.45,    283.45,  283.45,  283.45,
  283.45,    283.45,  283.45,  283.45,
  283.35,    283.35,  283.35,  283.35,
  283.3,     283.3,   283.3,   283.3,
  283.3,     283.3,   283.3,   283.3,
  283.3,     283.3,   283.3,   283.3,
  283.55,    283.55,  283.55,  283.55,
  283.85,    283.85,  283.85,  283.85,
  284.05,    284.05,  284.05,  284.05,
  284.2,     284.2,   284.2,   284.2,
  284.35,    284.35,  284.35,  284.35,
  284.3,     284.3,   284.3,   284.3,
  283.9,     283.9,   283.9,   283.9,
  283.65,    283.65,  283.65,  283.65,
  283.65,    283.65,  283.65,  283.65,
  283.6,     283.6,   283.6,   283.6,
  283.5,     283.5,   283.5,   283.5,
  283.35,    283.35,  283.35,  283.35,
  283,       283,     283,     283,
  282.25,    282.25,  282.25,  282.25,
  280.65,    280.65,  280.65,  280.65,
  279.35,    279.35,  279.35,  279.35,
  279.05,    279.05,  279.05,  279.05,
  278.65,    278.65,  278.65,  278.65,
  278.3,     278.3,   278.3,   278.3,
  278.35,    278.35,  278.35,  278.35,
  277.8,     277.8,   277.8,   277.8,
  277.8,     277.8,   277.8,   277.8,
  277.55,    277.55,  277.55,  277.55,
  276.9,     276.9,   276.9,   276.9,
  277.1,     277.1,   277.1,   277.1,
  277.25,    277.25,  277.25,  277.25,
  277.95,    277.95,  277.95,  277.95,
  279.6,     279.6,   279.6,   279.6,
  281.5,     281.5,   281.5,   281.5,
  282.1,     282.1,   282.1,   282.1,
  281.75,    281.75,  281.75,  281.75,
  281.55,    281.55,  281.55,  281.55,
  281.65,    281.65,  281.65,  281.65,
  282.15,    282.15,  282.15,  282.15,
  283.15,    283.15,  283.15,  283.15,
  284.2,     284.2,   284.2,   284.2,
  285,       285,     285,     285,
  285.85,    285.85,  285.85,  285.85,
  286.9,     286.9,   286.9,   286.9,
  287.5,     287.5,   287.5,   287.5,
  287.75,    287.75,  287.75,  287.75,
  288.4,     288.4,   288.4,   288.4,
  289.1,     289.1,   289.1,   289.1,
  289.55,    289.55,  289.55,  289.55,
  289.75,    289.75,  289.75,  289.75,
  290,       290,     290,     290,
  290.65,    290.65,  290.65,  290.65,
  291.1,     291.1,   291.1,   291.1,
  291.2,     291.2,   291.2,   291.2,
  291.2,     291.2,   291.2,   291.2,
  291.1,     291.1,   291.1,   291.1,
  290.9,     290.9,   290.9,   290.9,
  290.5,     290.5,   290.5,   290.5,
  289.95,    289.95,  289.95,  289.95,
  289.35,    289.35,  289.35,  289.35,
  288.7,     288.7,   288.7,   288.7,
  288.1,     288.1,   288.1,   288.1,
  287.65,    287.65,  287.65,  287.65,
  287.25,    287.25,  287.25,  287.25,
  286.95,    286.95,  286.95,  286.95,
  286.8,     286.8,   286.8,   286.8,
  286.65,    286.65,  286.65,  286.65,
  286.45,    286.45,  286.45,  286.45,
  286.3,     286.3,   286.3,   286.3,
  286.15,    286.15,  286.15,  286.15,
  285.95,    285.95,  285.95,  285.95,
  285.9,     285.9,   285.9,   285.9,
  286,       286,     286,     286,
  286,       286,     286,     286,
  285.95,    285.95,  285.95,  285.95,
  285.95,    285.95,  285.95,  285.95,
  286,       286,     286,     286,
  286.05,    286.05,  286.05,  286.05,
  286.15,    286.15,  286.15,  286.15,
  286.35,    286.35,  286.35,  286.35,
  286.6,     286.6,   286.6,   286.6,
  287.05,    287.05,  287.05,  287.05,
  287.85,    287.85,  287.85,  287.85,
  288.65,    288.65,  288.65,  288.65,
  289.4,     289.4,   289.4,   289.4,
  290.15,    290.15,  290.15,  290.15,
  290.95,    290.95,  290.95,  290.95,
  292.1,     292.1,   292.1,   292.1,
  293,       293,     293,     293,
  293.7,     293.7,   293.7,   293.7,
  294.5,     294.5,   294.5,   294.5,
  295.05,    295.05,  295.05,  295.05,
  295.6,     295.6,   295.6,   295.6,
  296.15,    296.15,  296.15,  296.15,
  296.55,    296.55,  296.55,  296.55,
  296.65,    296.65,  296.65,  296.65,
  296.6,     296.6,   296.6,   296.6,
  296.95,    296.95,  296.95,  296.95,
  297.45,    297.45,  297.45,  297.45,
  297.7,     297.7,   297.7,   297.7,
  297.8,     297.8,   297.8,   297.8,
  297.9,     297.9,   297.9,   297.9,
  297.85,    297.85,  297.85,  297.85,
  297.6,     297.6,   297.6,   297.6,
  297.25,    297.25,  297.25,  297.25,
  296.8,     296.8,   296.8,   296.8,
  296.35,    296.35,  296.35,  296.35,
  295.85,    295.85,  295.85,  295.85,
  295.25,    295.25,  295.25,  295.25,
  294.55,    294.55,  294.55,  294.55,
  293.9,     293.9,   293.9,   293.9,
  293.3,     293.3,   293.3,   293.3,
  292.75,    292.75,  292.75,  292.75,
  292.35,    292.35,  292.35,  292.35,
  292.25,    292.25,  292.25,  292.25,
  292.05,    292.05,  292.05,  292.05,
  291.55,    291.55,  291.55,  291.55,
  291.25,    291.25,  291.25,  291.25,
  290.85,    290.85,  290.85,  290.85,
  290.5,     290.5,   290.5,   290.5,
  290.25,    290.25,  290.25,  290.25,
  290.05,    290.05,  290.05,  290.05,
  290.3,     290.3,   290.3,   290.3,
  290,       290,     290,     290,
  289.3,     289.3,   289.3,   289.3,
  289,       289,     289,     289,
  288.9,     288.9,   288.9,   288.9,
  289.25,    289.25,  289.25,  289.25,
  289.9,     289.9,   289.9,   289.9,
  290.7,     290.7,   290.7,   290.7,
  291.7,     291.7,   291.7,   291.7,
  292.9,     292.9,   292.9,   292.9,
  293.8,     293.8,   293.8,   293.8,
  294.25,    294.25,  294.25,  294.25,
  294.7,     294.7,   294.7,   294.7,
  295.3,     295.3,   295.3,   295.3,
  296,       296,     296,     296,
  296.55,    296.55,  296.55,  296.55,
  297.2,     297.2,   297.2,   297.2,
  298,       298,     298,     298,
  298.5,     298.5,   298.5,   298.5,
  298.9,     298.9,   298.9,   298.9,
  299.4,     299.4,   299.4,   299.4,
  299.85,    299.85,  299.85,  299.85,
  300.15,    300.15,  300.15,  300.15,
  300.35,    300.35,  300.35,  300.35,
  300.4,     300.4,   300.4,   300.4,
  300.45,    300.45,  300.45,  300.45,
  300.65,    300.65,  300.65,  300.65,
  300.75,    300.75,  300.75,  300.75,
  300.75,    300.75,  300.75,  300.75,
  300.75,    300.75,  300.75,  300.75,
  300.8,     300.8,   300.8,   300.8,
  299.95,    299.95,  299.95,  299.95,
  298.05,    298.05,  298.05,  298.05,
  296.7,     296.7,   296.7,   296.7,
  296.35,    296.35,  296.35,  296.35,
  296.3,     296.3,   296.3,   296.3,
  295.55,    295.55,  295.55,  295.55,
  294.7,     294.7,   294.7,   294.7,
  295.05,    295.05,  295.05,  295.05,
  295.15,    295.15,  295.15,  295.15,
  294.65,    294.65,  294.65,  294.65,
  294.05,    294.05,  294.05,  294.05,
  292.55,    292.55,  292.55,  292.55,
  292,       292,     292,     292,
  292.65,    292.65,  292.65,  292.65,
  292.2,     292.2,   292.2,   292.2,
  291.9,     291.9,   291.9,   291.9,
  291.85,    291.85,  291.85,  291.85,
  291.3,     291.3,   291.3,   291.3,
  290.85,    290.85,  290.85,  290.85,
  290.25,    290.25,  290.25,  290.25,
  289.8,     289.8,   289.8,   289.8,
  289.65,    289.65,  289.65,  289.65,
  289.6,     289.6,   289.6,   289.6,
  289.8,     289.8,   289.8,   289.8,
  290.3,     290.3,   290.3,   290.3,
  290.95,    290.95,  290.95,  290.95,
  291.55,    291.55,  291.55,  291.55,
  291.95,    291.95,  291.95,  291.95,
  292.45,    292.45,  292.45,  292.45,
  293.15,    293.15,  293.15,  293.15,
  293.35,    293.35,  293.35,  293.35,
  293.1,     293.1,   293.1,   293.1,
  293.2,     293.2,   293.2,   293.2,
  293.45,    293.45,  293.45,  293.45,
  293.35,    293.35,  293.35,  293.35,
  292.95,    292.95,  292.95,  292.95,
  292.6,     292.6,   292.6,   292.6,
  292.15,    292.15,  292.15,  292.15,
  291.7,     291.7,   291.7,   291.7,
  290.65,    290.65,  290.65,  290.65,
  289.45,    289.45,  289.45,  289.45,
  289.3,     289.3,   289.3,   289.3,
  289.55,    289.55,  289.55,  289.55,
  289.8,     289.8,   289.8,   289.8,
  290.05,    290.05,  290.05,  290.05,
  290.3,     290.3,   290.3,   290.3,
  290.4,     290.4,   290.4,   290.4,
  290.4,     290.4,   290.4,   290.4,
  290.3,     290.3,   290.3,   290.3,
  290.15,    290.15,  290.15,  290.15,
  290.15,    290.15,  290.15,  290.15,
  290,       290,     290,     290,
  289.6,     289.6,   289.6,   289.6,
  289.1,     289.1,   289.1,   289.1,
  288.65,    288.65,  288.65,  288.65,
  288.4,     288.4,   288.4,   288.4,
  288.35,    288.35,  288.35,  288.35,
  288.25,    288.25,  288.25,  288.25,
  288.05,    288.05,  288.05,  288.05,
  287.9,     287.9,   287.9,   287.9,
  287.9,     287.9,   287.9,   287.9,
  288.05,    288.05,  288.05,  288.05,
  288.3,     288.3,   288.3,   288.3,
  288.5,     288.5,   288.5,   288.5,
  288.45,    288.45,  288.45,  288.45,
  288.25,    288.25,  288.25,  288.25,
  288.1,     288.1,   288.1,   288.1,
  287.9,     287.9,   287.9,   287.9,
  287.65,    287.65,  287.65,  287.65,
  287.45,    287.45,  287.45,  287.45,
  287.4,     287.4,   287.4,   287.4,
  287.5,     287.5,   287.5,   287.5,
  287.6,     287.6,   287.6,   287.6,
  287.9,     287.9,   287.9,   287.9,
  288.25,    288.25,  288.25,  288.25,
  288.6,     288.6,   288.6,   288.6,
  288.8,     288.8,   288.8,   288.8,
  289.05,    289.05,  289.05,  289.05,
  289.65,    289.65,  289.65,  289.65,
  290.35,    290.35,  290.35,  290.35,
  290.95,    290.95,  290.95,  290.95,
  291.3,     291.3,   291.3,   291.3,
  291.9,     291.9,   291.9,   291.9,
  292.4,     292.4,   292.4,   292.4,
  292.65,    292.65,  292.65,  292.65,
  293.1,     293.1,   293.1,   293.1,
  293.65,    293.65,  293.65,  293.65,
  294.25,    294.25,  294.25,  294.25,
  294.6,     294.6,   294.6,   294.6,
  294.55,    294.55,  294.55,  294.55,
  294.75,    294.75,  294.75,  294.75,
  295.15,    295.15,  295.15,  295.15,
  295.3,     295.3,   295.3,   295.3,
  295.35,    295.35,  295.35,  295.35,
  295.1,     295.1,   295.1,   295.1,
  294.8,     294.8,   294.8,   294.8,
  294.6,     294.6,   294.6,   294.6,
  294.2,     294.2,   294.2,   294.2,
  293.45,    293.45,  293.45,  293.45,
  291.75,    291.75,  291.75,  291.75,
  289.4,     289.4,   289.4,   289.4,
  288.1,     288.1,   288.1,   288.1,
  287.85,    287.85,  287.85,  287.85,
  287.65,    287.65,  287.65,  287.65,
  287.55,    287.55,  287.55,  287.55,
  287.55,    287.55,  287.55,  287.55,
  287.55,    287.55,  287.55,  287.55,
  287.55,    287.55,  287.55,  287.55,
  287.45,    287.45,  287.45,  287.45,
  287.25,    287.25,  287.25,  287.25,
  287,       287,     287,     287,
  286.95,    286.95,  286.95,  286.95,
  287.15,    287.15,  287.15,  287.15,
  287.25,    287.25,  287.25,  287.25,
  287.15,    287.15,  287.15,  287.15,
  286.95,    286.95,  286.95,  286.95,
  286.85,    286.85,  286.85,  286.85,
  286.8,     286.8,   286.8,   286.8,
  286.75,    286.75,  286.75,  286.75,
  286.9,     286.9,   286.9,   286.9,
  287.25,    287.25,  287.25,  287.25,
  287.55,    287.55,  287.55,  287.55,
  287.95,    287.95,  287.95,  287.95,
  288.65,    288.65,  288.65,  288.65,
  289.05,    289.05,  289.05,  289.05,
  289.15,    289.15,  289.15,  289.15,
  289.45,    289.45,  289.45,  289.45,
  289.8,     289.8,   289.8,   289.8,
  290.1,     290.1,   290.1,   290.1,
  290.95,    290.95,  290.95,  290.95,
  291.9,     291.9,   291.9,   291.9,
  292.45,    292.45,  292.45,  292.45,
  292.85,    292.85,  292.85,  292.85,
  292.8,     292.8,   292.8,   292.8,
  291.95,    291.95,  291.95,  291.95,
  289.3,     289.3,   289.3,   289.3,
  287.2,     287.2,   287.2,   287.2,
  287.4,     287.4,   287.4,   287.4,
  287.85,    287.85,  287.85,  287.85,
  287.8,     287.8,   287.8,   287.8,
  287.45,    287.45,  287.45,  287.45,
  287.2,     287.2,   287.2,   287.2,
  287.2,     287.2,   287.2,   287.2,
  287.35,    287.35,  287.35,  287.35,
  287.35,    287.35,  287.35,  287.35,
  287,       287,     287,     287,
  286.5,     286.5,   286.5,   286.5,
  285.6,     285.6,   285.6,   285.6,
  284.8,     284.8,   284.8,   284.8,
  284.5,     284.5,   284.5,   284.5,
  284.2,     284.2,   284.2,   284.2,
  283.9,     283.9,   283.9,   283.9,
  283.55,    283.55,  283.55,  283.55,
  283.35,    283.35,  283.35,  283.35,
  283.3,     283.3,   283.3,   283.3,
  283.2,     283.2,   283.2,   283.2,
  283.35,    283.35,  283.35,  283.35,
  283.9,     283.9,   283.9,   283.9,
  284.4,     284.4,   284.4,   284.4,
  284.55,    284.55,  284.55,  284.55,
  284.55,    284.55,  284.55,  284.55,
  284.5,     284.5,   284.5,   284.5,
  284.3,     284.3,   284.3,   284.3,
  284.05,    284.05,  284.05,  284.05,
  284.1,     284.1,   284.1,   284.1,
  284.5,     284.5,   284.5,   284.5,
  284.7,     284.7,   284.7,   284.7,
  284.6,     284.6,   284.6,   284.6,
  284.5,     284.5,   284.5,   284.5,
  284.5,     284.5,   284.5,   284.5,
  284.6,     284.6,   284.6,   284.6,
  284.75,    284.75,  284.75,  284.75,
  284.8,     284.8,   284.8,   284.8,
  284.75,    284.75,  284.75,  284.75,
  284.85,    284.85,  284.85,  284.85,
  285,       285,     285,     285,
  285.2,     285.2,   285.2,   285.2,
  285.45,    285.45,  285.45,  285.45,
  285.8,     285.8,   285.8,   285.8,
  286.25,    286.25,  286.25,  286.25,
  286.95,    286.95,  286.95,  286.95,
  287.95,    287.95,  287.95,  287.95,
  288.5,     288.5,   288.5,   288.5,
  287.8,     287.8,   287.8,   287.8,
  286.65,    286.65,  286.65,  286.65,
  286.45,    286.45,  286.45,  286.45,
  286.4,     286.4,   286.4,   286.4,
  285.85,    285.85,  285.85,  285.85,
  285.3,     285.3,   285.3,   285.3,
  285.1,     285.1,   285.1,   285.1,
  285.1,     285.1,   285.1,   285.1,
  284.8,     284.8,   284.8,   284.8,
  284.35,    284.35,  284.35,  284.35,
  283.9,     283.9,   283.9,   283.9,
  283.35,    283.35,  283.35,  283.35,
  282.9,     282.9,   282.9,   282.9,
  282.65,    282.65,  282.65,  282.65,
  282.5,     282.5,   282.5,   282.5,
  282.4,     282.4,   282.4,   282.4,
  282.25,    282.25,  282.25,  282.25,
  282.1,     282.1,   282.1,   282.1,
  281.95,    281.95,  281.95,  281.95,
  281.8,     281.8,   281.8,   281.8,
  281.75,    281.75,  281.75,  281.75,
  281.8,     281.8,   281.8,   281.8,
  281.9,     281.9,   281.9,   281.9,
  282,       282,     282,     282,
  282.1,     282.1,   282.1,   282.1,
  282.2,     282.2,   282.2,   282.2,
  282.25,    282.25,  282.25,  282.25,
  282.25,    282.25,  282.25,  282.25,
  282.25,    282.25,  282.25,  282.25,
  282.3,     282.3,   282.3,   282.3,
  282.4,     282.4,   282.4,   282.4,
  282.6,     282.6,   282.6,   282.6,
  282.9,     282.9,   282.9,   282.9,
  283.2,     283.2,   283.2,   283.2,
  283.5,     283.5,   283.5,   283.5,
  283.7,     283.7,   283.7,   283.7,
  283.9,     283.9,   283.9,   283.9,
  284.3,     284.3,   284.3,   284.3,
  284.4,     284.4,   284.4,   284.4,
  284.3,     284.3,   284.3,   284.3,
  284.3,     284.3,   284.3,   284.3,
  284.25,    284.25,  284.25,  284.25,
  284.2,     284.2,   284.2,   284.2,
  284.3,     284.3,   284.3,   284.3,
  284.5,     284.5,   284.5,   284.5,
  284.65,    284.65,  284.65,  284.65,
  284.7,     284.7,   284.7,   284.7,
  284.55,    284.55,  284.55,  284.55,
  284.35,    284.35,  284.35,  284.35,
  284.55,    284.55,  284.55,  284.55,
  284.9,     284.9,   284.9,   284.9,
  284.85,    284.85,  284.85,  284.85,
  284.8,     284.8,   284.8,   284.8,
  284.8,     284.8,   284.8,   284.8,
  284.4,     284.4,   284.4,   284.4,
  284,       284,     284,     284,
  284,       284,     284,     284,
  283.8,     283.8,   283.8,   283.8,
  283.5,     283.5,   283.5,   283.5,
  283.3,     283.3,   283.3,   283.3,
  282.95,    282.95,  282.95,  282.95,
  282.55,    282.55,  282.55,  282.55,
  282.2,     282.2,   282.2,   282.2,
  281.95,    281.95,  281.95,  281.95,
  281.75,    281.75,  281.75,  281.75,
  281.45,    281.45,  281.45,  281.45,
  281.1,     281.1,   281.1,   281.1,
  280.95,    280.95,  280.95,  280.95,
  280.85,    280.85,  280.85,  280.85,
  280.8,     280.8,   280.8,   280.8,
  280.7,     280.7,   280.7,   280.7,
  280.45,    280.45,  280.45,  280.45,
  280.25,    280.25,  280.25,  280.25,
  280.05,    280.05,  280.05,  280.05,
  279.65,    279.65,  279.65,  279.65,
  279.3,     279.3,   279.3,   279.3,
  279.25,    279.25,  279.25,  279.25,
  279,       279,     279,     279,
  278.85,    278.85,  278.85,  278.85,
  279.35,    279.35,  279.35,  279.35,
  280.4,     280.4,   280.4,   280.4,
  281.7,     281.7,   281.7,   281.7,
  282.65,    282.65,  282.65,  282.65,
  283.1,     283.1,   283.1,   283.1,
  283.2,     283.2,   283.2,   283.2,
  283.1,     283.1,   283.1,   283.1,
  283.2,     283.2,   283.2,   283.2,
  283.65,    283.65,  283.65,  283.65,
  284.1,     284.1,   284.1,   284.1,
  284.05,    284.05,  284.05,  284.05,
  284.3,     284.3,   284.3,   284.3,
  284.75,    284.75,  284.75,  284.75,
  284.95,    284.95,  284.95,  284.95,
  285.45,    285.45,  285.45,  285.45,
  285.45,    285.45,  285.45,  285.45,
  285.45,    285.45,  285.45,  285.45,
  285.5,     285.5,   285.5,   285.5,
  285.45,    285.45,  285.45,  285.45,
  285.45,    285.45,  285.45,  285.45,
  285.35,    285.35,  285.35,  285.35,
  285.55,    285.55,  285.55,  285.55,
  285.45,    285.45,  285.45,  285.45,
  285.2,     285.2,   285.2,   285.2,
  285,       285,     285,     285,
  284.6,     284.6,   284.6,   284.6,
  284.15,    284.15,  284.15,  284.15,
  283.65,    283.65,  283.65,  283.65,
  282.9,     282.9,   282.9,   282.9,
  282,       282,     282,     282,
  281.1,     281.1,   281.1,   281.1,
  280.45,    280.45,  280.45,  280.45,
  280,       280,     280,     280,
  279.6,     279.6,   279.6,   279.6,
  279.15,    279.15,  279.15,  279.15,
  278.6,     278.6,   278.6,   278.6,
  278.3,     278.3,   278.3,   278.3,
  278.15,    278.15,  278.15,  278.15,
  278.1,     278.1,   278.1,   278.1,
  278.1,     278.1,   278.1,   278.1,
  277.95,    277.95,  277.95,  277.95,
  277.5,     277.5,   277.5,   277.5,
  276.9,     276.9,   276.9,   276.9,
  276.9,     276.9,   276.9,   276.9,
  277.1,     277.1,   277.1,   277.1,
  277.05,    277.05,  277.05,  277.05,
  277.35,    277.35,  277.35,  277.35,
  278.1,     278.1,   278.1,   278.1,
  279.25,    279.25,  279.25,  279.25,
  280.25,    280.25,  280.25,  280.25,
  280.9,     280.9,   280.9,   280.9,
  281.4,     281.4,   281.4,   281.4,
  281.9,     281.9,   281.9,   281.9,
  282.25,    282.25,  282.25,  282.25,
  282.5,     282.5,   282.5,   282.5,
  282.75,    282.75,  282.75,  282.75,
  282.95,    282.95,  282.95,  282.95,
  283.3,     283.3,   283.3,   283.3,
  283.7,     283.7,   283.7,   283.7,
  283.95,    283.95,  283.95,  283.95,
  284.2,     284.2,   284.2,   284.2,
  284.7,     284.7,   284.7,   284.7,
  285.3,     285.3,   285.3,   285.3,
  285.65,    285.65,  285.65,  285.65,
  285.95,    285.95,  285.95,  285.95,
  286.3,     286.3,   286.3,   286.3,
  286.35,    286.35,  286.35,  286.35,
  286.45,    286.45,  286.45,  286.45,
  286.7,     286.7,   286.7,   286.7,
  286.9,     286.9,   286.9,   286.9,
  286.95,    286.95,  286.95,  286.95,
  286.75,    286.75,  286.75,  286.75,
  286.7,     286.7,   286.7,   286.7,
  286.7,     286.7,   286.7,   286.7,
  286.3,     286.3,   286.3,   286.3,
  285.95,    285.95,  285.95,  285.95,
  285.55,    285.55,  285.55,  285.55,
  284.95,    284.95,  284.95,  284.95,
  284.1,     284.1,   284.1,   284.1,
  283.05,    283.05,  283.05,  283.05,
  282,       282,     282,     282,
  281.15,    281.15,  281.15,  281.15,
  280.65,    280.65,  280.65,  280.65,
  280.25,    280.25,  280.25,  280.25,
  279.95,    279.95,  279.95,  279.95,
  280.2,     280.2,   280.2,   280.2,
  280.55,    280.55,  280.55,  280.55,
  280.4,     280.4,   280.4,   280.4,
  280.05,    280.05,  280.05,  280.05,
  279.7,     279.7,   279.7,   279.7,
  279.5,     279.5,   279.5,   279.5,
  279.4,     279.4,   279.4,   279.4,
  279.2,     279.2,   279.2,   279.2,
  278.9,     278.9,   278.9,   278.9,
  278.75,    278.75,  278.75,  278.75,
  279.15,    279.15,  279.15,  279.15,
  280.15,    280.15,  280.15,  280.15,
  281.55,    281.55,  281.55,  281.55,
  283.3,     283.3,   283.3,   283.3,
  284.8,     284.8,   284.8,   284.8,
  285.65,    285.65,  285.65,  285.65,
  286.35,    286.35,  286.35,  286.35,
  286.85,    286.85,  286.85,  286.85,
  287.05,    287.05,  287.05,  287.05,
  287.15,    287.15,  287.15,  287.15,
  287.1,     287.1,   287.1,   287.1,
  287.25,    287.25,  287.25,  287.25,
  287.6,     287.6,   287.6,   287.6,
  287.95,    287.95,  287.95,  287.95,
  288.2,     288.2,   288.2,   288.2,
  288.45,    288.45,  288.45,  288.45,
  288.75,    288.75,  288.75,  288.75,
  289.15,    289.15,  289.15,  289.15,
  289.55,    289.55,  289.55,  289.55,
  289.65,    289.65,  289.65,  289.65,
  289.7,     289.7,   289.7,   289.7,
  289.95,    289.95,  289.95,  289.95,
  290,       290,     290,     290,
  289.75,    289.75,  289.75,  289.75,
  289.65,    289.65,  289.65,  289.65,
  289.45,    289.45,  289.45,  289.45,
  289.25,    289.25,  289.25,  289.25,
  288.85,    288.85,  288.85,  288.85,
  287.75,    287.75,  287.75,  287.75,
  286.65,    286.65,  286.65,  286.65,
  285.85,    285.85,  285.85,  285.85,
  285.05,    285.05,  285.05,  285.05,
  284.25,    284.25,  284.25,  284.25,
  283.45,    283.45,  283.45,  283.45,
  282.7,     282.7,   282.7,   282.7,
  282.05,    282.05,  282.05,  282.05,
  281.5,     281.5,   281.5,   281.5,
  281.05,    281.05,  281.05,  281.05,
  280.55,    280.55,  280.55,  280.55,
  279.85,    279.85,  279.85,  279.85,
  279.2,     279.2,   279.2,   279.2,
  278.7,     278.7,   278.7,   278.7,
  278.45,    278.45,  278.45,  278.45,
  278.25,    278.25,  278.25,  278.25,
  278.15,    278.15,  278.15,  278.15,
  278.1,     278.1,   278.1,   278.1,
  277.85,    277.85,  277.85,  277.85,
  278.1,     278.1,   278.1,   278.1,
  278.05,    278.05,  278.05,  278.05,
  278,       278,     278,     278,
  279.15,    279.15,  279.15,  279.15,
  280.65,    280.65,  280.65,  280.65,
  281.7,     281.7,   281.7,   281.7,
  282.55,    282.55,  282.55,  282.55,
  283.35,    283.35,  283.35,  283.35,
  284.05,    284.05,  284.05,  284.05,
  284.6,     284.6,   284.6,   284.6,
  284.95,    284.95,  284.95,  284.95,
  285.25,    285.25,  285.25,  285.25,
  285.55,    285.55,  285.55,  285.55,
  286,       286,     286,     286,
  286.65,    286.65,  286.65,  286.65,
  287.3,     287.3,   287.3,   287.3,
  287.85,    287.85,  287.85,  287.85,
  288.2,     288.2,   288.2,   288.2,
  288.4,     288.4,   288.4,   288.4,
  288.7,     288.7,   288.7,   288.7,
  288.95,    288.95,  288.95,  288.95,
  289.1,     289.1,   289.1,   289.1,
  289.1,     289.1,   289.1,   289.1,
  288.95,    288.95,  288.95,  288.95,
  288.65,    288.65,  288.65,  288.65,
  288.35,    288.35,  288.35,  288.35,
  288.15,    288.15,  288.15,  288.15,
  287.95,    287.95,  287.95,  287.95,
  287.65,    287.65,  287.65,  287.65,
  287.2,     287.2,   287.2,   287.2,
  286.7,     286.7,   286.7,   286.7,
  286.2,     286.2,   286.2,   286.2,
  285.8,     285.8,   285.8,   285.8,
  285.55,    285.55,  285.55,  285.55,
  285.3,     285.3,   285.3,   285.3,
  285,       285,     285,     285,
  284.7,     284.7,   284.7,   284.7,
  284.45,    284.45,  284.45,  284.45,
  284.4,     284.4,   284.4,   284.4,
  284.35,    284.35,  284.35,  284.35,
  284.05,    284.05,  284.05,  284.05,
  283.65,    283.65,  283.65,  283.65,
  283.35,    283.35,  283.35,  283.35,
  283.15,    283.15,  283.15,  283.15,
  283,       283,     283,     283,
  282.95,    282.95,  282.95,  282.95,
  282.9,     282.9,   282.9,   282.9,
  282.9,     282.9,   282.9,   282.9,
  282.95,    282.95,  282.95,  282.95,
  282.85,    282.85,  282.85,  282.85,
  282.7,     282.7,   282.7,   282.7,
  282.45,    282.45,  282.45,  282.45,
  282.35,    282.35,  282.35,  282.35,
  282.5,     282.5,   282.5,   282.5,
  282.65,    282.65,  282.65,  282.65,
  282.85,    282.85,  282.85,  282.85,
  283.05,    283.05,  283.05,  283.05,
  283.45,    283.45,  283.45,  283.45,
  283.7,     283.7,   283.7,   283.7,
  283.65,    283.65,  283.65,  283.65,
  283.75,    283.75,  283.75,  283.75,
  283.95,    283.95,  283.95,  283.95,
  284.1,     284.1,   284.1,   284.1,
  284.2,     284.2,   284.2,   284.2,
  284.1,     284.1,   284.1,   284.1,
  284.05,    284.05,  284.05,  284.05,
  284.25,    284.25,  284.25,  284.25,
  284.25,    284.25,  284.25,  284.25,
  284.05,    284.05,  284.05,  284.05,
  284,       284,     284,     284,
  284.25,    284.25,  284.25,  284.25,
  284.45,    284.45,  284.45,  284.45,
  284.35,    284.35,  284.35,  284.35,
  284.15,    284.15,  284.15,  284.15,
  284,       284,     284,     284,
  283.8,     283.8,   283.8,   283.8,
  283.55,    283.55,  283.55,  283.55,
  283.3,     283.3,   283.3,   283.3,
  283.05,    283.05,  283.05,  283.05,
  282.8,     282.8,   282.8,   282.8,
  282.55,    282.55,  282.55,  282.55,
  282.45,    282.45,  282.45,  282.45,
  282.35,    282.35,  282.35,  282.35,
  282.2,     282.2,   282.2,   282.2,
  282.05,    282.05,  282.05,  282.05,
  281.9,     281.9,   281.9,   281.9,
  281.95,    281.95,  281.95,  281.95,
  282,       282,     282,     282,
  281.9,     281.9,   281.9,   281.9,
  281.8,     281.8,   281.8,   281.8,
  281.65,    281.65,  281.65,  281.65,
  281.5,     281.5,   281.5,   281.5,
  281.45,    281.45,  281.45,  281.45,
  281.5,     281.5,   281.5,   281.5,
  281.45,    281.45,  281.45,  281.45,
  281.15,    281.15,  281.15,  281.15,
  280.95,    280.95,  280.95,  280.95,
  281.05,    281.05,  281.05,  281.05,
  281.4,     281.4,   281.4,   281.4,
  281.8,     281.8,   281.8,   281.8,
  282.05,    282.05,  282.05,  282.05,
  282.25,    282.25,  282.25,  282.25,
  282.7,     282.7,   282.7,   282.7,
  283.4,     283.4,   283.4,   283.4,
  284.05,    284.05,  284.05,  284.05,
  284.35,    284.35,  284.35,  284.35,
  284.35,    284.35,  284.35,  284.35,
  284.65,    284.65,  284.65,  284.65,
  285.05,    285.05,  285.05,  285.05,
  285.35,    285.35,  285.35,  285.35,
  285.75,    285.75,  285.75,  285.75,
  286.1,     286.1,   286.1,   286.1,
  286.4,     286.4,   286.4,   286.4,
  286.55,    286.55,  286.55,  286.55,
  286.6,     286.6,   286.6,   286.6,
  286.8,     286.8,   286.8,   286.8,
  286.9,     286.9,   286.9,   286.9,
  286.9,     286.9,   286.9,   286.9,
  287,       287,     287,     287,
  287.1,     287.1,   287.1,   287.1,
  287.2,     287.2,   287.2,   287.2,
  287.35,    287.35,  287.35,  287.35,
  287.4,     287.4,   287.4,   287.4,
  287.15,    287.15,  287.15,  287.15,
  286.75,    286.75,  286.75,  286.75,
  286.1,     286.1,   286.1,   286.1,
  285.2,     285.2,   285.2,   285.2,
  284.3,     284.3,   284.3,   284.3,
  283.45,    283.45,  283.45,  283.45,
  282.7,     282.7,   282.7,   282.7,
  282.05,    282.05,  282.05,  282.05,
  281.45,    281.45,  281.45,  281.45,
  280.95,    280.95,  280.95,  280.95,
  280.5,     280.5,   280.5,   280.5,
  280.15,    280.15,  280.15,  280.15,
  279.9,     279.9,   279.9,   279.9,
  279.6,     279.6,   279.6,   279.6,
  279.3,     279.3,   279.3,   279.3,
  279,       279,     279,     279,
  278.7,     278.7,   278.7,   278.7,
  278.35,    278.35,  278.35,  278.35,
  278.1,     278.1,   278.1,   278.1,
  278,       278,     278,     278,
  277.7,     277.7,   277.7,   277.7,
  277.85,    277.85,  277.85,  277.85,
  278.45,    278.45,  278.45,  278.45,
  278.95,    278.95,  278.95,  278.95,
  279.9,     279.9,   279.9,   279.9,
  281.15,    281.15,  281.15,  281.15,
  282.05,    282.05,  282.05,  282.05,
  282.55,    282.55,  282.55,  282.55,
  282.9,     282.9,   282.9,   282.9,
  283.3,     283.3,   283.3,   283.3,
  283.8,     283.8,   283.8,   283.8,
  284.3,     284.3,   284.3,   284.3,
  285.05,    285.05,  285.05,  285.05,
  285.85,    285.85,  285.85,  285.85,
  286.4,     286.4,   286.4,   286.4,
  286.95,    286.95,  286.95,  286.95,
  287.4,     287.4,   287.4,   287.4,
  288,       288,     288,     288,
  288.7,     288.7,   288.7,   288.7,
  288.95,    288.95,  288.95,  288.95,
  288.95,    288.95,  288.95,  288.95,
  289.05,    289.05,  289.05,  289.05,
  289.45,    289.45,  289.45,  289.45,
  289.7,     289.7,   289.7,   289.7,
  289.45,    289.45,  289.45,  289.45,
  288.9,     288.9,   288.9,   288.9,
  288.25,    288.25,  288.25,  288.25,
  287.9,     287.9,   287.9,   287.9,
  287.9,     287.9,   287.9,   287.9,
  287.65,    287.65,  287.65,  287.65,
  286.85,    286.85,  286.85,  286.85,
  285.85,    285.85,  285.85,  285.85,
  285.05,    285.05,  285.05,  285.05,
  284.45,    284.45,  284.45,  284.45,
  283.85,    283.85,  283.85,  283.85,
  283.35,    283.35,  283.35,  283.35,
  282.95,    282.95,  282.95,  282.95,
  282.6,     282.6,   282.6,   282.6,
  282.3,     282.3,   282.3,   282.3,
  281.95,    281.95,  281.95,  281.95,
  281.6,     281.6,   281.6,   281.6,
  281.35,    281.35,  281.35,  281.35,
  281.3,     281.3,   281.3,   281.3,
  281.4,     281.4,   281.4,   281.4,
  281.5,     281.5,   281.5,   281.5,
  281.5,     281.5,   281.5,   281.5,
  281.5,     281.5,   281.5,   281.5,
  281.5,     281.5,   281.5,   281.5,
  281.35,    281.35,  281.35,  281.35,
  281.35,    281.35,  281.35,  281.35,
  281.6,     281.6,   281.6,   281.6,
  281.85,    281.85,  281.85,  281.85,
  282.05,    282.05,  282.05,  282.05,
  282.1,     282.1,   282.1,   282.1,
  282.3,     282.3,   282.3,   282.3,
  282.95,    282.95,  282.95,  282.95,
  283.85,    283.85,  283.85,  283.85,
  284.65,    284.65,  284.65,  284.65,
  285.6,     285.6,   285.6,   285.6,
  286.85,    286.85,  286.85,  286.85,
  287.75,    287.75,  287.75,  287.75,
  288.35,    288.35,  288.35,  288.35,
  288.95,    288.95,  288.95,  288.95,
  289.5,     289.5,   289.5,   289.5,
  290.2,     290.2,   290.2,   290.2,
  290.65,    290.65,  290.65,  290.65,
  290.9,     290.9,   290.9,   290.9,
  291.35,    291.35,  291.35,  291.35,
  291.7,     291.7,   291.7,   291.7,
  291.95,    291.95,  291.95,  291.95,
  292.15,    292.15,  292.15,  292.15,
  292.35,    292.35,  292.35,  292.35,
  292.4,     292.4,   292.4,   292.4,
  292.3,     292.3,   292.3,   292.3,
  292.25,    292.25,  292.25,  292.25,
  292.15,    292.15,  292.15,  292.15,
  291.95,    291.95,  291.95,  291.95,
  291.7,     291.7,   291.7,   291.7,
  291.3,     291.3,   291.3,   291.3,
  290.65,    290.65,  290.65,  290.65,
  289.75,    289.75,  289.75,  289.75,
  288.75,    288.75,  288.75,  288.75,
  287.75,    287.75,  287.75,  287.75,
  286.65,    286.65,  286.65,  286.65,
  285.9,     285.9,   285.9,   285.9,
  285.6,     285.6,   285.6,   285.6,
  285.1,     285.1,   285.1,   285.1,
  284.55,    284.55,  284.55,  284.55,
  284,       284,     284,     284,
  283.55,    283.55,  283.55,  283.55,
  283.3,     283.3,   283.3,   283.3,
  283,       283,     283,     283,
  282.7,     282.7,   282.7,   282.7,
  282.4,     282.4,   282.4,   282.4,
  282.15,    282.15,  282.15,  282.15,
  281.85,    281.85,  281.85,  281.85,
  281.6,     281.6,   281.6,   281.6,
  281.55,    281.55,  281.55,  281.55,
  281.7,     281.7,   281.7,   281.7,
  282.35,    282.35,  282.35,  282.35,
  283.1,     283.1,   283.1,   283.1,
  283.8,     283.8,   283.8,   283.8,
  285.3,     285.3,   285.3,   285.3,
  286.7,     286.7,   286.7,   286.7,
  287.3,     287.3,   287.3,   287.3,
  287.65,    287.65,  287.65,  287.65,
  287.9,     287.9,   287.9,   287.9,
  288.15,    288.15,  288.15,  288.15,
  288.45,    288.45,  288.45,  288.45,
  288.8,     288.8,   288.8,   288.8,
  289.1,     289.1,   289.1,   289.1,
  289.35,    289.35,  289.35,  289.35,
  289.55,    289.55,  289.55,  289.55,
  289.8,     289.8,   289.8,   289.8,
  289.85,    289.85,  289.85,  289.85,
  289.95,    289.95,  289.95,  289.95,
  290.1,     290.1,   290.1,   290.1,
  290.15,    290.15,  290.15,  290.15,
  290.3,     290.3,   290.3,   290.3,
  290.45,    290.45,  290.45,  290.45,
  290.5,     290.5,   290.5,   290.5,
  290.45,    290.45,  290.45,  290.45,
  290.25,    290.25,  290.25,  290.25,
  289.9,     289.9,   289.9,   289.9,
  289.65,    289.65,  289.65,  289.65,
  289.45,    289.45,  289.45,  289.45,
  289.2,     289.2,   289.2,   289.2,
  288.65,    288.65,  288.65,  288.65,
  287.75,    287.75,  287.75,  287.75,
  286.8,     286.8,   286.8,   286.8,
  286,       286,     286,     286,
  285.8,     285.8,   285.8,   285.8,
  286,       286,     286,     286,
  285.8,     285.8,   285.8,   285.8,
  285.25,    285.25,  285.25,  285.25,
  284.6,     284.6,   284.6,   284.6,
  283.9,     283.9,   283.9,   283.9,
  283.2,     283.2,   283.2,   283.2,
  282.65,    282.65,  282.65,  282.65,
  282.3,     282.3,   282.3,   282.3,
  281.9,     281.9,   281.9,   281.9,
  281.4,     281.4,   281.4,   281.4,
  280.95,    280.95,  280.95,  280.95,
  280.6,     280.6,   280.6,   280.6,
  280.5,     280.5,   280.5,   280.5,
  280.65,    280.65,  280.65,  280.65,
  280.9,     280.9,   280.9,   280.9,
  281.3,     281.3,   281.3,   281.3,
  281.9,     281.9,   281.9,   281.9,
  282.65,    282.65,  282.65,  282.65,
  283.4,     283.4,   283.4,   283.4,
  284.15,    284.15,  284.15,  284.15,
  285,       285,     285,     285,
  285.85,    285.85,  285.85,  285.85,
  286.5,     286.5,   286.5,   286.5,
  287.2,     287.2,   287.2,   287.2,
  287.85,    287.85,  287.85,  287.85,
  288.3,     288.3,   288.3,   288.3,
  288.9,     288.9,   288.9,   288.9,
  289.55,    289.55,  289.55,  289.55,
  290.05,    290.05,  290.05,  290.05,
  290.4,     290.4,   290.4,   290.4,
  290.8,     290.8,   290.8,   290.8,
  291.3,     291.3,   291.3,   291.3,
  291.75,    291.75,  291.75,  291.75,
  291.85,    291.85,  291.85,  291.85,
  291.9,     291.9,   291.9,   291.9,
  292.1,     292.1,   292.1,   292.1,
  292.2,     292.2,   292.2,   292.2,
  292.25,    292.25,  292.25,  292.25,
  292.25,    292.25,  292.25,  292.25,
  292.15,    292.15,  292.15,  292.15,
  291.8,     291.8,   291.8,   291.8,
  291.45,    291.45,  291.45,  291.45,
  290.7,     290.7,   290.7,   290.7,
  289.85,    289.85,  289.85,  289.85,
  289.5,     289.5,   289.5,   289.5,
  289.1,     289.1,   289.1,   289.1,
  288.6,     288.6,   288.6,   288.6,
  288.3,     288.3,   288.3,   288.3,
  288.25,    288.25,  288.25,  288.25,
  288.1,     288.1,   288.1,   288.1,
  287.75,    287.75,  287.75,  287.75,
  287.3,     287.3,   287.3,   287.3,
  286.9,     286.9,   286.9,   286.9,
  286.6,     286.6,   286.6,   286.6,
  286.15,    286.15,  286.15,  286.15,
  285.65,    285.65,  285.65,  285.65,
  285.3,     285.3,   285.3,   285.3,
  285.05,    285.05,  285.05,  285.05,
  284.75,    284.75,  284.75,  284.75,
  284.35,    284.35,  284.35,  284.35,
  284,       284,     284,     284,
  283.8,     283.8,   283.8,   283.8,
  283.85,    283.85,  283.85,  283.85,
  284.2,     284.2,   284.2,   284.2,
  284.7,     284.7,   284.7,   284.7,
  285.25,    285.25,  285.25,  285.25,
  285.95,    285.95,  285.95,  285.95,
  286.7,     286.7,   286.7,   286.7,
  287.6,     287.6,   287.6,   287.6,
  288.6,     288.6,   288.6,   288.6,
  289.45,    289.45,  289.45,  289.45,
  290.05,    290.05,  290.05,  290.05,
  290.55,    290.55,  290.55,  290.55,
  291.15,    291.15,  291.15,  291.15,
  291.65,    291.65,  291.65,  291.65,
  291.95,    291.95,  291.95,  291.95,
  292.15,    292.15,  292.15,  292.15,
  292.35,    292.35,  292.35,  292.35,
  292.55,    292.55,  292.55,  292.55,
  292.75,    292.75,  292.75,  292.75,
  293.05,    293.05,  293.05,  293.05,
  293.25,    293.25,  293.25,  293.25,
  293.35,    293.35,  293.35,  293.35,
  293.5,     293.5,   293.5,   293.5,
  293.55,    293.55,  293.55,  293.55,
  293.6,     293.6,   293.6,   293.6,
  293.7,     293.7,   293.7,   293.7,
  293.65,    293.65,  293.65,  293.65,
  293.55,    293.55,  293.55,  293.55,
  293.35,    293.35,  293.35,  293.35,
  292.9,     292.9,   292.9,   292.9,
  292.15,    292.15,  292.15,  292.15,
  291.05,    291.05,  291.05,  291.05,
  290.05,    290.05,  290.05,  290.05,
  289.2,     289.2,   289.2,   289.2,
  288.35,    288.35,  288.35,  288.35,
  287.4,     287.4,   287.4,   287.4,
  286.75,    286.75,  286.75,  286.75,
  286.75,    286.75,  286.75,  286.75,
  286.7,     286.7,   286.7,   286.7,
  286.3,     286.3,   286.3,   286.3,
  285.8,     285.8,   285.8,   285.8,
  285.4,     285.4,   285.4,   285.4,
  285,       285,     285,     285,
  284.65,    284.65,  284.65,  284.65,
  284.25,    284.25,  284.25,  284.25,
  283.7,     283.7,   283.7,   283.7,
  283.05,    283.05,  283.05,  283.05,
  282.4,     282.4,   282.4,   282.4,
  282.05,    282.05,  282.05,  282.05,
  282.35,    282.35,  282.35,  282.35,
  283.6,     283.6,   283.6,   283.6,
  285.3,     285.3,   285.3,   285.3,
  286.8,     286.8,   286.8,   286.8,
  287.9,     287.9,   287.9,   287.9,
  289.1,     289.1,   289.1,   289.1,
  290.15,    290.15,  290.15,  290.15,
  290.75,    290.75,  290.75,  290.75,
  291.25,    291.25,  291.25,  291.25,
  291.7,     291.7,   291.7,   291.7,
  292.1,     292.1,   292.1,   292.1,
  292.55,    292.55,  292.55,  292.55,
  293,       293,     293,     293,
  293.25,    293.25,  293.25,  293.25,
  293.55,    293.55,  293.55,  293.55,
  293.8,     293.8,   293.8,   293.8,
  294.1,     294.1,   294.1,   294.1,
  294.3,     294.3,   294.3,   294.3,
  294.4,     294.4,   294.4,   294.4,
  294.55,    294.55,  294.55,  294.55,
  294.75,    294.75,  294.75,  294.75,
  294.9,     294.9,   294.9,   294.9,
  294.85,    294.85,  294.85,  294.85,
  294.9,     294.9,   294.9,   294.9,
  294.95,    294.95,  294.95,  294.95,
  294.8,     294.8,   294.8,   294.8,
  294.45,    294.45,  294.45,  294.45,
  294.25,    294.25,  294.25,  294.25,
  294.05,    294.05,  294.05,  294.05,
  293.45,    293.45,  293.45,  293.45,
  292,       292,     292,     292,
  290.2,     290.2,   290.2,   290.2,
  289.1,     289.1,   289.1,   289.1,
  288.4,     288.4,   288.4,   288.4,
  287.75,    287.75,  287.75,  287.75,
  287.2,     287.2,   287.2,   287.2,
  286.65,    286.65,  286.65,  286.65,
  286.15,    286.15,  286.15,  286.15,
  285.9,     285.9,   285.9,   285.9,
  285.75,    285.75,  285.75,  285.75,
  285.5,     285.5,   285.5,   285.5,
  285.15,    285.15,  285.15,  285.15,
  284.75,    284.75,  284.75,  284.75,
  284.4,     284.4,   284.4,   284.4,
  284.25,    284.25,  284.25,  284.25,
  284.35,    284.35,  284.35,  284.35,
  283.7,     283.7,   283.7,   283.7,
  282.45,    282.45,  282.45,  282.45,
  282.15,    282.15,  282.15,  282.15,
  282.85,    282.85,  282.85,  282.85,
  284.05,    284.05,  284.05,  284.05,
  285.4,     285.4,   285.4,   285.4,
  286.75,    286.75,  286.75,  286.75,
  288.1,     288.1,   288.1,   288.1,
  289.2,     289.2,   289.2,   289.2,
  290.3,     290.3,   290.3,   290.3,
  291.35,    291.35,  291.35,  291.35,
  292.4,     292.4,   292.4,   292.4,
  293.25,    293.25,  293.25,  293.25,
  293.5,     293.5,   293.5,   293.5,
  293.6,     293.6,   293.6,   293.6,
  293.75,    293.75,  293.75,  293.75,
  294,       294,     294,     294,
  294.2,     294.2,   294.2,   294.2,
  294.5,     294.5,   294.5,   294.5,
  294.8,     294.8,   294.8,   294.8,
  294.65,    294.65,  294.65,  294.65,
  294.7,     294.7,   294.7,   294.7,
  295.05,    295.05,  295.05,  295.05,
  295.25,    295.25,  295.25,  295.25,
  295.2,     295.2,   295.2,   295.2,
  295.05,    295.05,  295.05,  295.05,
  295.15,    295.15,  295.15,  295.15,
  295.1,     295.1,   295.1,   295.1,
  294.5,     294.5,   294.5,   294.5,
  293.75,    293.75,  293.75,  293.75,
  293.1,     293.1,   293.1,   293.1,
  292.25,    292.25,  292.25,  292.25,
  291.25,    291.25,  291.25,  291.25,
  290.1,     290.1,   290.1,   290.1,
  289.2,     289.2,   289.2,   289.2,
  288.75,    288.75,  288.75,  288.75,
  288.3,     288.3,   288.3,   288.3,
  287.9,     287.9,   287.9,   287.9,
  287.6,     287.6,   287.6,   287.6,
  287.3,     287.3,   287.3,   287.3,
  287,       287,     287,     287,
  286.65,    286.65,  286.65,  286.65,
  286.35,    286.35,  286.35,  286.35,
  286.25,    286.25,  286.25,  286.25,
  286.1,     286.1,   286.1,   286.1,
  285.85,    285.85,  285.85,  285.85,
  285.65,    285.65,  285.65,  285.65,
  285.45,    285.45,  285.45,  285.45,
  285.45,    285.45,  285.45,  285.45,
  285.7,     285.7,   285.7,   285.7,
  286.15,    286.15,  286.15,  286.15,
  286.55,    286.55,  286.55,  286.55,
  287.05,    287.05,  287.05,  287.05,
  288.1,     288.1,   288.1,   288.1,
  289.55,    289.55,  289.55,  289.55,
  291.6,     291.6,   291.6,   291.6,
  293.5,     293.5,   293.5,   293.5,
  294.7,     294.7,   294.7,   294.7,
  295.6,     295.6,   295.6,   295.6,
  296.15,    296.15,  296.15,  296.15,
  296.55,    296.55,  296.55,  296.55,
  296.7,     296.7,   296.7,   296.7,
  297.05,    297.05,  297.05,  297.05,
  297.55,    297.55,  297.55,  297.55,
  297.9,     297.9,   297.9,   297.9,
  298.3,     298.3,   298.3,   298.3,
  298.55,    298.55,  298.55,  298.55,
  298.6,     298.6,   298.6,   298.6,
  298.65,    298.65,  298.65,  298.65,
  298.85,    298.85,  298.85,  298.85,
  298.85,    298.85,  298.85,  298.85,
  298.85,    298.85,  298.85,  298.85,
  298.85,    298.85,  298.85,  298.85,
  298.65,    298.65,  298.65,  298.65,
  298.5,     298.5,   298.5,   298.5,
  298.2,     298.2,   298.2,   298.2,
  297.8,     297.8,   297.8,   297.8,
  297.45,    297.45,  297.45,  297.45,
  296.9,     296.9,   296.9,   296.9,
  296.2,     296.2,   296.2,   296.2,
  295.45,    295.45,  295.45,  295.45,
  294.8,     294.8,   294.8,   294.8,
  294.35,    294.35,  294.35,  294.35,
  293.95,    293.95,  293.95,  293.95,
  293.75,    293.75,  293.75,  293.75,
  293.6,     293.6,   293.6,   293.6,
  293.2,     293.2,   293.2,   293.2,
  292.65,    292.65,  292.65,  292.65,
  292,       292,     292,     292,
  291.35,    291.35,  291.35,  291.35,
  290.8,     290.8,   290.8,   290.8,
  290.3,     290.3,   290.3,   290.3,
  289.9,     289.9,   289.9,   289.9,
  289.55,    289.55,  289.55,  289.55,
  289.2,     289.2,   289.2,   289.2,
  288.9,     288.9,   288.9,   288.9,
  288.65,    288.65,  288.65,  288.65,
  288.65,    288.65,  288.65,  288.65,
  289.2,     289.2,   289.2,   289.2,
  290,       290,     290,     290,
  290.4,     290.4,   290.4,   290.4,
  290.85,    290.85,  290.85,  290.85,
  291.65,    291.65,  291.65,  291.65,
  292.4,     292.4,   292.4,   292.4,
  292.85,    292.85,  292.85,  292.85,
  293.3,     293.3,   293.3,   293.3,
  294,       294,     294,     294,
  295,       295,     295,     295,
  296.2,     296.2,   296.2,   296.2,
  297.1,     297.1,   297.1,   297.1,
  297.8,     297.8,   297.8,   297.8,
  298.3,     298.3,   298.3,   298.3,
  298.75,    298.75,  298.75,  298.75,
  299.25,    299.25,  299.25,  299.25,
  299.55,    299.55,  299.55,  299.55,
  299.85,    299.85,  299.85,  299.85,
  300,       300,     300,     300,
  299.8,     299.8,   299.8,   299.8,
  299.95,    299.95,  299.95,  299.95,
  300.25,    300.25,  300.25,  300.25,
  299.95,    299.95,  299.95,  299.95,
  299.65,    299.65,  299.65,  299.65,
  299.55,    299.55,  299.55,  299.55,
  299.5,     299.5,   299.5,   299.5,
  299.55,    299.55,  299.55,  299.55,
  299.45,    299.45,  299.45,  299.45,
  299.15,    299.15,  299.15,  299.15,
  298.5,     298.5,   298.5,   298.5,
  297.65,    297.65,  297.65,  297.65,
  296.85,    296.85,  296.85,  296.85,
  296.15,    296.15,  296.15,  296.15,
  295.2,     295.2,   295.2,   295.2,
  294.75,    294.75,  294.75,  294.75,
  295.05,    295.05,  295.05,  295.05,
  295,       295,     295,     295,
  294.7,     294.7,   294.7,   294.7,
  294.5,     294.5,   294.5,   294.5,
  294.2,     294.2,   294.2,   294.2,
  293.7,     293.7,   293.7,   293.7,
  293.35,    293.35,  293.35,  293.35,
  293.2,     293.2,   293.2,   293.2,
  293.1,     293.1,   293.1,   293.1,
  292.85,    292.85,  292.85,  292.85,
  292.45,    292.45,  292.45,  292.45,
  292.05,    292.05,  292.05,  292.05,
  291.9,     291.9,   291.9,   291.9,
  292.2,     292.2,   292.2,   292.2,
  292.5,     292.5,   292.5,   292.5,
  292.65,    292.65,  292.65,  292.65,
  293.3,     293.3,   293.3,   293.3,
  294.35,    294.35,  294.35,  294.35,
  295.25,    295.25,  295.25,  295.25,
  296.05,    296.05,  296.05,  296.05,
  296.8,     296.8,   296.8,   296.8,
  297.45,    297.45,  297.45,  297.45,
  298.2,     298.2,   298.2,   298.2,
  298.9,     298.9,   298.9,   298.9,
  299.3,     299.3,   299.3,   299.3,
  299.75,    299.75,  299.75,  299.75,
  300,       300,     300,     300,
  300.2,     300.2,   300.2,   300.2,
  300.7,     300.7,   300.7,   300.7,
  301.2,     301.2,   301.2,   301.2,
  301.2,     301.2,   301.2,   301.2,
  300.95,    300.95,  300.95,  300.95,
  300.75,    300.75,  300.75,  300.75,
  296.65,    296.65,  296.65,  296.65,
  291.45,    291.45,  291.45,  291.45,
  290.1,     290.1,   290.1,   290.1,
  290.45,    290.45,  290.45,  290.45,
  291.3,     291.3,   291.3,   291.3,
  291.8,     291.8,   291.8,   291.8,
  291.9,     291.9,   291.9,   291.9,
  292,       292,     292,     292,
  291.95,    291.95,  291.95,  291.95,
  291.9,     291.9,   291.9,   291.9,
  291.8,     291.8,   291.8,   291.8,
  291.85,    291.85,  291.85,  291.85,
  291.85,    291.85,  291.85,  291.85,
  291.45,    291.45,  291.45,  291.45,
  290.9,     290.9,   290.9,   290.9,
  290.55,    290.55,  290.55,  290.55,
  290.2,     290.2,   290.2,   290.2,
  290,       290,     290,     290,
  290,       290,     290,     290,
  289.85,    289.85,  289.85,  289.85,
  289.8,     289.8,   289.8,   289.8,
  289.7,     289.7,   289.7,   289.7,
  289.5,     289.5,   289.5,   289.5,
  289.45,    289.45,  289.45,  289.45,
  289.65,    289.65,  289.65,  289.65,
  289.75,    289.75,  289.75,  289.75,
  289.7,     289.7,   289.7,   289.7,
  289.75,    289.75,  289.75,  289.75,
  289.85,    289.85,  289.85,  289.85,
  289.85,    289.85,  289.85,  289.85,
  289.85,    289.85,  289.85,  289.85,
  289.8,     289.8,   289.8,   289.8,
  289.9,     289.9,   289.9,   289.9,
  290.1,     290.1,   290.1,   290.1,
  290.25,    290.25,  290.25,  290.25,
  290.4,     290.4,   290.4,   290.4,
  290.45,    290.45,  290.45,  290.45,
  290.35,    290.35,  290.35,  290.35,
  290.35,    290.35,  290.35,  290.35,
  290.55,    290.55,  290.55,  290.55,
  290.8,     290.8,   290.8,   290.8,
  291.05,    291.05,  291.05,  291.05,
  290.85,    290.85,  290.85,  290.85,
  290,       290,     290,     290,
  289.7,     289.7,   289.7,   289.7,
  289.95,    289.95,  289.95,  289.95,
  290.1,     290.1,   290.1,   290.1,
  290.5,     290.5,   290.5,   290.5,
  291,       291,     291,     291,
  291.5,     291.5,   291.5,   291.5,
  291.9,     291.9,   291.9,   291.9,
  292.25,    292.25,  292.25,  292.25,
  292.7,     292.7,   292.7,   292.7,
  292.8,     292.8,   292.8,   292.8,
  292.25,    292.25,  292.25,  292.25,
  291.85,    291.85,  291.85,  291.85,
  291.75,    291.75,  291.75,  291.75,
  291.55,    291.55,  291.55,  291.55,
  291.05,    291.05,  291.05,  291.05,
  290.3,     290.3,   290.3,   290.3,
  289.65,    289.65,  289.65,  289.65,
  289.25,    289.25,  289.25,  289.25,
  289,       289,     289,     289,
  288.5,     288.5,   288.5,   288.5,
  287.75,    287.75,  287.75,  287.75,
  286.95,    286.95,  286.95,  286.95,
  286.25,    286.25,  286.25,  286.25,
  285.75,    285.75,  285.75,  285.75,
  285.5,     285.5,   285.5,   285.5,
  285.35,    285.35,  285.35,  285.35,
  284.95,    284.95,  284.95,  284.95,
  284.6,     284.6,   284.6,   284.6,
  284.5,     284.5,   284.5,   284.5,
  284.4,     284.4,   284.4,   284.4,
  284.45,    284.45,  284.45,  284.45,
  284.7,     284.7,   284.7,   284.7,
  285.15,    285.15,  285.15,  285.15,
  285.85,    285.85,  285.85,  285.85,
  286.5,     286.5,   286.5,   286.5,
  286.95,    286.95,  286.95,  286.95,
  287.45,    287.45,  287.45,  287.45,
  288.05,    288.05,  288.05,  288.05,
  288.6,     288.6,   288.6,   288.6,
  288.8,     288.8,   288.8,   288.8,
  289.05,    289.05,  289.05,  289.05,
  289.9,     289.9,   289.9,   289.9,
  290.65,    290.65,  290.65,  290.65,
  291.3,     291.3,   291.3,   291.3,
  291.75,    291.75,  291.75,  291.75,
  291.9,     291.9,   291.9,   291.9,
  292.35,    292.35,  292.35,  292.35,
  292.8,     292.8,   292.8,   292.8,
  293.15,    293.15,  293.15,  293.15,
  293.35,    293.35,  293.35,  293.35,
  293.6,     293.6,   293.6,   293.6,
  293.9,     293.9,   293.9,   293.9,
  294,       294,     294,     294,
  293.9,     293.9,   293.9,   293.9,
  293.7,     293.7,   293.7,   293.7,
  293.8,     293.8,   293.8,   293.8,
  293.85,    293.85,  293.85,  293.85,
  293.75,    293.75,  293.75,  293.75,
  293.7,     293.7,   293.7,   293.7,
  293.45,    293.45,  293.45,  293.45,
  292.65,    292.65,  292.65,  292.65,
  291.6,     291.6,   291.6,   291.6,
  290.65,    290.65,  290.65,  290.65,
  289.6,     289.6,   289.6,   289.6,
  288.7,     288.7,   288.7,   288.7,
  287.9,     287.9,   287.9,   287.9,
  287.15,    287.15,  287.15,  287.15,
  286.7,     286.7,   286.7,   286.7,
  286.4,     286.4,   286.4,   286.4,
  286.05,    286.05,  286.05,  286.05,
  285.9,     285.9,   285.9,   285.9,
  286,       286,     286,     286,
  285.95,    285.95,  285.95,  285.95,
  285.8,     285.8,   285.8,   285.8,
  285.65,    285.65,  285.65,  285.65,
  285.5,     285.5,   285.5,   285.5,
  285.35,    285.35,  285.35,  285.35,
  285.15,    285.15,  285.15,  285.15,
  285.05,    285.05,  285.05,  285.05,
  285.05,    285.05,  285.05,  285.05,
  285.3,     285.3,   285.3,   285.3,
  286,       286,     286,     286,
  287.05,    287.05,  287.05,  287.05,
  288.1,     288.1,   288.1,   288.1,
  288.95,    288.95,  288.95,  288.95,
  289.75,    289.75,  289.75,  289.75,
  290.65,    290.65,  290.65,  290.65,
  291.65,    291.65,  291.65,  291.65,
  292.45,    292.45,  292.45,  292.45,
  293,       293,     293,     293,
  293.55,    293.55,  293.55,  293.55,
  294.05,    294.05,  294.05,  294.05,
  294.5,     294.5,   294.5,   294.5,
  294.9,     294.9,   294.9,   294.9,
  295.3,     295.3,   295.3,   295.3,
  295.75,    295.75,  295.75,  295.75,
  296,       296,     296,     296,
  296.1,     296.1,   296.1,   296.1,
  296.35,    296.35,  296.35,  296.35,
  296.6,     296.6,   296.6,   296.6,
  296.8,     296.8,   296.8,   296.8,
  297,       297,     297,     297,
  297.1,     297.1,   297.1,   297.1,
  297.15,    297.15,  297.15,  297.15,
  297.2,     297.2,   297.2,   297.2,
  297.1,     297.1,   297.1,   297.1,
  296.8,     296.8,   296.8,   296.8,
  296.45,    296.45,  296.45,  296.45,
  296.05,    296.05,  296.05,  296.05,
  295.5,     295.5,   295.5,   295.5,
  294.95,    294.95,  294.95,  294.95,
  294.55,    294.55,  294.55,  294.55,
  294.05,    294.05,  294.05,  294.05,
  293.4,     293.4,   293.4,   293.4,
  292.75,    292.75,  292.75,  292.75,
  292.2,     292.2,   292.2,   292.2,
  291.85,    291.85,  291.85,  291.85,
  291.7,     291.7,   291.7,   291.7,
  291.6,     291.6,   291.6,   291.6,
  291.4,     291.4,   291.4,   291.4,
  291.15,    291.15,  291.15,  291.15,
  290.9,     290.9,   290.9,   290.9,
  290.55,    290.55,  290.55,  290.55,
  290.25,    290.25,  290.25,  290.25,
  290.1,     290.1,   290.1,   290.1,
  290.05,    290.05,  290.05,  290.05,
  289.95,    289.95,  289.95,  289.95,
  289.95,    289.95,  289.95,  289.95,
  290.25,    290.25,  290.25,  290.25,
  290.55,    290.55,  290.55,  290.55,
  291,       291,     291,     291,
  291.5,     291.5,   291.5,   291.5,
  291.85,    291.85,  291.85,  291.85,
  292.25,    292.25,  292.25,  292.25,
  292.6,     292.6,   292.6,   292.6,
  292.85,    292.85,  292.85,  292.85,
  293.55,    293.55,  293.55,  293.55,
  294.65,    294.65,  294.65,  294.65,
  295.55,    295.55,  295.55,  295.55,
  296.3,     296.3,   296.3,   296.3,
  296.75,    296.75,  296.75,  296.75,
  296.9,     296.9,   296.9,   296.9,
  297,       297,     297,     297,
  297.1,     297.1,   297.1,   297.1,
  297.2,     297.2,   297.2,   297.2,
  297.35,    297.35,  297.35,  297.35,
  296.8,     296.8,   296.8,   296.8,
  294.15,    294.15,  294.15,  294.15,
  292.25,    292.25,  292.25,  292.25,
  292.5,     292.5,   292.5,   292.5,
  292.5,     292.5,   292.5,   292.5,
  292.25,    292.25,  292.25,  292.25,
  292.1,     292.1,   292.1,   292.1,
  292,       292,     292,     292,
  291.9,     291.9,   291.9,   291.9,
  291.85,    291.85,  291.85,  291.85,
  291.8,     291.8,   291.8,   291.8,
  291.7,     291.7,   291.7,   291.7,
  291.55,    291.55,  291.55,  291.55,
  291.35,    291.35,  291.35,  291.35,
  291.25,    291.25,  291.25,  291.25,
  291.15,    291.15,  291.15,  291.15,
  291.1,     291.1,   291.1,   291.1,
  291.15,    291.15,  291.15,  291.15,
  291.1,     291.1,   291.1,   291.1,
  291.1,     291.1,   291.1,   291.1,
  291.05,    291.05,  291.05,  291.05,
  290.2,     290.2,   290.2,   290.2,
  289.1,     289.1,   289.1,   289.1,
  288.5,     288.5,   288.5,   288.5,
  288.15,    288.15,  288.15,  288.15,
  288,       288,     288,     288,
  287.95,    287.95,  287.95,  287.95,
  288.05,    288.05,  288.05,  288.05,
  288.2,     288.2,   288.2,   288.2,
  288.2,     288.2,   288.2,   288.2,
  288.15,    288.15,  288.15,  288.15,
  288.2,     288.2,   288.2,   288.2,
  288.25,    288.25,  288.25,  288.25,
  288.4,     288.4,   288.4,   288.4,
  288.65,    288.65,  288.65,  288.65,
  289.15,    289.15,  289.15,  289.15,
  289.85,    289.85,  289.85,  289.85,
  290.25,    290.25,  290.25,  290.25,
  290.45,    290.45,  290.45,  290.45,
  290.95,    290.95,  290.95,  290.95,
  291.6,     291.6,   291.6,   291.6,
  292.2,     292.2,   292.2,   292.2,
  292.7,     292.7,   292.7,   292.7,
  293.05,    293.05,  293.05,  293.05,
  293.5,     293.5,   293.5,   293.5,
  293.5,     293.5,   293.5,   293.5,
  292.9,     292.9,   292.9,   292.9,
  292.55,    292.55,  292.55,  292.55,
  292.95,    292.95,  292.95,  292.95,
  293.7,     293.7,   293.7,   293.7,
  293.45,    293.45,  293.45,  293.45,
  292.85,    292.85,  292.85,  292.85,
  292.9,     292.9,   292.9,   292.9,
  292.9,     292.9,   292.9,   292.9,
  292.9,     292.9,   292.9,   292.9,
  292.85,    292.85,  292.85,  292.85,
  292.75,    292.75,  292.75,  292.75,
  292.9,     292.9,   292.9,   292.9,
  292.9,     292.9,   292.9,   292.9,
  292.45,    292.45,  292.45,  292.45,
  291.9,     291.9,   291.9,   291.9,
  291.45,    291.45,  291.45,  291.45,
  291.1,     291.1,   291.1,   291.1,
  290.75,    290.75,  290.75,  290.75,
  290.4,     290.4,   290.4,   290.4,
  290.1,     290.1,   290.1,   290.1,
  289.75,    289.75,  289.75,  289.75,
  289.45,    289.45,  289.45,  289.45,
  289.25,    289.25,  289.25,  289.25,
  288.95,    288.95,  288.95,  288.95,
  288.65,    288.65,  288.65,  288.65,
  288.4,     288.4,   288.4,   288.4,
  288.25,    288.25,  288.25,  288.25,
  288.2,     288.2,   288.2,   288.2,
  288.05,    288.05,  288.05,  288.05,
  287.95,    287.95,  287.95,  287.95,
  287.95,    287.95,  287.95,  287.95,
  287.9,     287.9,   287.9,   287.9,
  287.9,     287.9,   287.9,   287.9,
  287.95,    287.95,  287.95,  287.95,
  288.05,    288.05,  288.05,  288.05,
  288.2,     288.2,   288.2,   288.2,
  288.55,    288.55,  288.55,  288.55,
  289.3,     289.3,   289.3,   289.3,
  289.9,     289.9,   289.9,   289.9,
  290.25,    290.25,  290.25,  290.25,
  290.95,    290.95,  290.95,  290.95,
  291.55,    291.55,  291.55,  291.55,
  291.95,    291.95,  291.95,  291.95,
  292.4,     292.4,   292.4,   292.4,
  292.5,     292.5,   292.5,   292.5,
  292.5,     292.5,   292.5,   292.5,
  292.9,     292.9,   292.9,   292.9,
  293.5,     293.5,   293.5,   293.5,
  293.9,     293.9,   293.9,   293.9,
  294.1,     294.1,   294.1,   294.1,
  294.05,    294.05,  294.05,  294.05,
  293.25,    293.25,  293.25,  293.25,
  292.9,     292.9,   292.9,   292.9,
  292.8,     292.8,   292.8,   292.8,
  291.5,     291.5,   291.5,   291.5,
  290.4,     290.4,   290.4,   290.4,
  290.4,     290.4,   290.4,   290.4,
  290.85,    290.85,  290.85,  290.85,
  290.95,    290.95,  290.95,  290.95,
  290.75,    290.75,  290.75,  290.75,
  290.6,     290.6,   290.6,   290.6,
  290.55,    290.55,  290.55,  290.55,
  290.55,    290.55,  290.55,  290.55,
  290.25,    290.25,  290.25,  290.25,
  289.8,     289.8,   289.8,   289.8,
  289.7,     289.7,   289.7,   289.7,
  289.55,    289.55,  289.55,  289.55,
  289.1,     289.1,   289.1,   289.1,
  288.7,     288.7,   288.7,   288.7,
  288.5,     288.5,   288.5,   288.5,
  288.35,    288.35,  288.35,  288.35,
  288.05,    288.05,  288.05,  288.05,
  287.8,     287.8,   287.8,   287.8,
  287.7,     287.7,   287.7,   287.7,
  287.7,     287.7,   287.7,   287.7,
  287.65,    287.65,  287.65,  287.65,
  287.45,    287.45,  287.45,  287.45,
  287.25,    287.25,  287.25,  287.25,
  287.15,    287.15,  287.15,  287.15,
  287.2,     287.2,   287.2,   287.2,
  287.3,     287.3,   287.3,   287.3,
  287.4,     287.4,   287.4,   287.4,
  287.45,    287.45,  287.45,  287.45,
  287.7,     287.7,   287.7,   287.7,
  288.1,     288.1,   288.1,   288.1,
  288.25,    288.25,  288.25,  288.25,
  288.35,    288.35,  288.35,  288.35,
  288.75,    288.75,  288.75,  288.75,
  289.05,    289.05,  289.05,  289.05,
  289.35,    289.35,  289.35,  289.35,
  289.75,    289.75,  289.75,  289.75,
  290.2,     290.2,   290.2,   290.2,
  290.75,    290.75,  290.75,  290.75,
  291.1,     291.1,   291.1,   291.1,
  291.45,    291.45,  291.45,  291.45,
  291.35,    291.35,  291.35,  291.35,
  290.4,     290.4,   290.4,   290.4,
  290.05,    290.05,  290.05,  290.05,
  290.2,     290.2,   290.2,   290.2,
  289.75,    289.75,  289.75,  289.75,
  288.95,    288.95,  288.95,  288.95,
  288.7,     288.7,   288.7,   288.7,
  288.85,    288.85,  288.85,  288.85,
  288.75,    288.75,  288.75,  288.75,
  288.85,    288.85,  288.85,  288.85,
  288.65,    288.65,  288.65,  288.65,
  288.15,    288.15,  288.15,  288.15,
  287.85,    287.85,  287.85,  287.85,
  287.75,    287.75,  287.75,  287.75,
  287.6,     287.6,   287.6,   287.6,
  287.2,     287.2,   287.2,   287.2,
  286.65,    286.65,  286.65,  286.65,
  286.2,     286.2,   286.2,   286.2,
  286,       286,     286,     286,
  285.95,    285.95,  285.95,  285.95,
  285.9,     285.9,   285.9,   285.9,
  285.85,    285.85,  285.85,  285.85,
  285.85,    285.85,  285.85,  285.85,
  285.8,     285.8,   285.8,   285.8,
  285.75,    285.75,  285.75,  285.75,
  285.65,    285.65,  285.65,  285.65,
  285.5,     285.5,   285.5,   285.5,
  285.4,     285.4,   285.4,   285.4,
  285.3,     285.3,   285.3,   285.3,
  285.2,     285.2,   285.2,   285.2,
  285.1,     285.1,   285.1,   285.1,
  285.05,    285.05,  285.05,  285.05,
  284.9,     284.9,   284.9,   284.9,
  284.75,    284.75,  284.75,  284.75,
  284.75,    284.75,  284.75,  284.75,
  284.85,    284.85,  284.85,  284.85,
  285.1,     285.1,   285.1,   285.1,
  285.45,    285.45,  285.45,  285.45,
  285.75,    285.75,  285.75,  285.75,
  286,       286,     286,     286,
  286.15,    286.15,  286.15,  286.15,
  286.05,    286.05,  286.05,  286.05,
  286.05,    286.05,  286.05,  286.05,
  286.2,     286.2,   286.2,   286.2,
  286.45,    286.45,  286.45,  286.45,
  286.9,     286.9,   286.9,   286.9,
  287.45,    287.45,  287.45,  287.45,
  287.7,     287.7,   287.7,   287.7,
  287.8,     287.8,   287.8,   287.8,
  288,       288,     288,     288,
  288.05,    288.05,  288.05,  288.05,
  288.2,     288.2,   288.2,   288.2,
  288.5,     288.5,   288.5,   288.5,
  288.6,     288.6,   288.6,   288.6,
  288.4,     288.4,   288.4,   288.4,
  288.3,     288.3,   288.3,   288.3,
  288.2,     288.2,   288.2,   288.2,
  287.8,     287.8,   287.8,   287.8,
  287.4,     287.4,   287.4,   287.4,
  287.3,     287.3,   287.3,   287.3,
  287.3,     287.3,   287.3,   287.3,
  286.95,    286.95,  286.95,  286.95,
  286.25,    286.25,  286.25,  286.25,
  285.5,     285.5,   285.5,   285.5,
  285,       285,     285,     285,
  284.6,     284.6,   284.6,   284.6,
  283.95,    283.95,  283.95,  283.95,
  283.3,     283.3,   283.3,   283.3,
  283.05,    283.05,  283.05,  283.05,
  282.85,    282.85,  282.85,  282.85,
  282.3,     282.3,   282.3,   282.3,
  282.1,     282.1,   282.1,   282.1,
  282.2,     282.2,   282.2,   282.2,
  282.1,     282.1,   282.1,   282.1,
  282.05,    282.05,  282.05,  282.05,
  282.1,     282.1,   282.1,   282.1,
  282.1,     282.1,   282.1,   282.1,
  282,       282,     282,     282,
  281.9,     281.9,   281.9,   281.9,
  282.1,     282.1,   282.1,   282.1,
  282.4,     282.4,   282.4,   282.4,
  282.15,    282.15,  282.15,  282.15,
  283,       283,     283,     283,
  285.05,    285.05,  285.05,  285.05,
  285.95,    285.95,  285.95,  285.95,
  286.1,     286.1,   286.1,   286.1,
  286.3,     286.3,   286.3,   286.3,
  286.3,     286.3,   286.3,   286.3,
  286.7,     286.7,   286.7,   286.7,
  287.35,    287.35,  287.35,  287.35,
  287.75,    287.75,  287.75,  287.75,
  288.05,    288.05,  288.05,  288.05,
  288.35,    288.35,  288.35,  288.35,
  288.85,    288.85,  288.85,  288.85,
  289.25,    289.25,  289.25,  289.25,
  289.3,     289.3,   289.3,   289.3,
  289.6,     289.6,   289.6,   289.6,
  289.85,    289.85,  289.85,  289.85,
  289.75,    289.75,  289.75,  289.75,
  289.75,    289.75,  289.75,  289.75,
  289.7,     289.7,   289.7,   289.7,
  289.75,    289.75,  289.75,  289.75,
  290,       290,     290,     290,
  290.05,    290.05,  290.05,  290.05,
  289.85,    289.85,  289.85,  289.85,
  289.65,    289.65,  289.65,  289.65,
  289.6,     289.6,   289.6,   289.6,
  289.5,     289.5,   289.5,   289.5,
  289.25,    289.25,  289.25,  289.25,
  288.9,     288.9,   288.9,   288.9,
  288.3,     288.3,   288.3,   288.3,
  287.5,     287.5,   287.5,   287.5,
  286.45,    286.45,  286.45,  286.45,
  285.5,     285.5,   285.5,   285.5,
  284.85,    284.85,  284.85,  284.85,
  284.2,     284.2,   284.2,   284.2,
  283.6,     283.6,   283.6,   283.6,
  283.15,    283.15,  283.15,  283.15,
  282.7,     282.7,   282.7,   282.7,
  282.3,     282.3,   282.3,   282.3,
  282.05,    282.05,  282.05,  282.05,
  281.8,     281.8,   281.8,   281.8,
  281.45,    281.45,  281.45,  281.45,
  281.05,    281.05,  281.05,  281.05,
  280.7,     280.7,   280.7,   280.7,
  280.4,     280.4,   280.4,   280.4,
  280.25,    280.25,  280.25,  280.25,
  280.35,    280.35,  280.35,  280.35,
  280.5,     280.5,   280.5,   280.5,
  280.9,     280.9,   280.9,   280.9,
  281.95,    281.95,  281.95,  281.95,
  283.3,     283.3,   283.3,   283.3,
  284.35,    284.35,  284.35,  284.35,
  285.1,     285.1,   285.1,   285.1,
  285.6,     285.6,   285.6,   285.6,
  286.05,    286.05,  286.05,  286.05,
  286.5,     286.5,   286.5,   286.5,
  286.7,     286.7,   286.7,   286.7,
  287.05,    287.05,  287.05,  287.05,
  287.35,    287.35,  287.35,  287.35,
  287.65,    287.65,  287.65,  287.65,
  288.2,     288.2,   288.2,   288.2,
  288.65,    288.65,  288.65,  288.65,
  288.9,     288.9,   288.9,   288.9,
  289.15,    289.15,  289.15,  289.15,
  289.45,    289.45,  289.45,  289.45,
  289.75,    289.75,  289.75,  289.75,
  289.8,     289.8,   289.8,   289.8,
  289.85,    289.85,  289.85,  289.85,
  289.95,    289.95,  289.95,  289.95,
  289.8,     289.8,   289.8,   289.8,
  289.85,    289.85,  289.85,  289.85,
  290.15,    290.15,  290.15,  290.15,
  290.2,     290.2,   290.2,   290.2,
  289.65,    289.65,  289.65,  289.65,
  289,       289,     289,     289,
  288.5,     288.5,   288.5,   288.5,
  288,       288,     288,     288,
  287.4,     287.4,   287.4,   287.4,
  286.65,    286.65,  286.65,  286.65,
  285.75,    285.75,  285.75,  285.75,
  284.9,     284.9,   284.9,   284.9,
  284.25,    284.25,  284.25,  284.25,
  283.6,     283.6,   283.6,   283.6,
  282.85,    282.85,  282.85,  282.85,
  282.4,     282.4,   282.4,   282.4,
  281.95,    281.95,  281.95,  281.95,
  281.55,    281.55,  281.55,  281.55,
  281.25,    281.25,  281.25,  281.25,
  280.75,    280.75,  280.75,  280.75,
  280.6,     280.6,   280.6,   280.6,
  280.55,    280.55,  280.55,  280.55,
  279.95,    279.95,  279.95,  279.95,
  279.1,     279.1,   279.1,   279.1,
  279,       279,     279,     279,
  279.4,     279.4,   279.4,   279.4,
  279.5,     279.5,   279.5,   279.5,
  279.5,     279.5,   279.5,   279.5,
  279.6,     279.6,   279.6,   279.6,
  280,       280,     280,     280,
  280.4,     280.4,   280.4,   280.4,
  281.15,    281.15,  281.15,  281.15,
  283.2,     283.2,   283.2,   283.2,
  285.05,    285.05,  285.05,  285.05,
  285.85,    285.85,  285.85,  285.85,
  286.2,     286.2,   286.2,   286.2,
  286.15,    286.15,  286.15,  286.15,
  286.3,     286.3,   286.3,   286.3,
  286.95,    286.95,  286.95,  286.95,
  287.25,    287.25,  287.25,  287.25,
  287.55,    287.55,  287.55,  287.55,
  288.25,    288.25,  288.25,  288.25,
  288.7,     288.7,   288.7,   288.7,
  289,       289,     289,     289,
  289.15,    289.15,  289.15,  289.15,
  289.45,    289.45,  289.45,  289.45,
  290,       290,     290,     290,
  290.5,     290.5,   290.5,   290.5,
  290.45,    290.45,  290.45,  290.45,
  290.3,     290.3,   290.3,   290.3,
  290.55,    290.55,  290.55,  290.55,
  290.65,    290.65,  290.65,  290.65,
  290.65,    290.65,  290.65,  290.65,
  290.6,     290.6,   290.6,   290.6,
  290.55,    290.55,  290.55,  290.55,
  290.25,    290.25,  290.25,  290.25,
  289.8,     289.8,   289.8,   289.8,
  289,       289,     289,     289,
  287.8,     287.8,   287.8,   287.8,
  286.7,     286.7,   286.7,   286.7,
  285.8,     285.8,   285.8,   285.8,
  285.15,    285.15,  285.15,  285.15,
  284.6,     284.6,   284.6,   284.6,
  284.15,    284.15,  284.15,  284.15,
  283.95,    283.95,  283.95,  283.95,
  283.85,    283.85,  283.85,  283.85,
  283.75,    283.75,  283.75,  283.75,
  283.7,     283.7,   283.7,   283.7,
  283.55,    283.55,  283.55,  283.55,
  283.35,    283.35,  283.35,  283.35,
  283.15,    283.15,  283.15,  283.15,
  282.95,    282.95,  282.95,  282.95,
  282.65,    282.65,  282.65,  282.65,
  282.3,     282.3,   282.3,   282.3,
  282.4,     282.4,   282.4,   282.4,
  282.95,    282.95,  282.95,  282.95,
  283.65,    283.65,  283.65,  283.65,
  284.9,     284.9,   284.9,   284.9,
  286.45,    286.45,  286.45,  286.45,
  287.7,     287.7,   287.7,   287.7,
  288.7,     288.7,   288.7,   288.7,
  289.45,    289.45,  289.45,  289.45,
  290,       290,     290,     290,
  290.55,    290.55,  290.55,  290.55,
  291.1,     291.1,   291.1,   291.1,
  291.6,     291.6,   291.6,   291.6,
  291.95,    291.95,  291.95,  291.95,
  292.15,    292.15,  292.15,  292.15,
  292.25,    292.25,  292.25,  292.25,
  292.45,    292.45,  292.45,  292.45,
  292.7,     292.7,   292.7,   292.7,
  292.8,     292.8,   292.8,   292.8,
  293.05,    293.05,  293.05,  293.05,
  293.4,     293.4,   293.4,   293.4,
  293.55,    293.55,  293.55,  293.55,
  293.45,    293.45,  293.45,  293.45,
  293.45,    293.45,  293.45,  293.45,
  293.5,     293.5,   293.5,   293.5,
  293.45,    293.45,  293.45,  293.45,
  293.4,     293.4,   293.4,   293.4,
  293.25,    293.25,  293.25,  293.25,
  293.05,    293.05,  293.05,  293.05,
  292.8,     292.8,   292.8,   292.8,
  292.5,     292.5,   292.5,   292.5,
  292.05,    292.05,  292.05,  292.05,
  291.4,     291.4,   291.4,   291.4,
  290.75,    290.75,  290.75,  290.75,
  290.3,     290.3,   290.3,   290.3,
  289.95,    289.95,  289.95,  289.95,
  289.4,     289.4,   289.4,   289.4,
  288.65,    288.65,  288.65,  288.65,
  288,       288,     288,     288,
  287.6,     287.6,   287.6,   287.6,
  287.3,     287.3,   287.3,   287.3,
  286.95,    286.95,  286.95,  286.95,
  286.55,    286.55,  286.55,  286.55,
  286.15,    286.15,  286.15,  286.15,
  285.8,     285.8,   285.8,   285.8,
  285.5,     285.5,   285.5,   285.5,
  285.05,    285.05,  285.05,  285.05,
  284.65,    284.65,  284.65,  284.65,
  284.55,    284.55,  284.55,  284.55,
  284.3,     284.3,   284.3,   284.3,
  283.9,     283.9,   283.9,   283.9,
  283.8,     283.8,   283.8,   283.8,
  283.85,    283.85,  283.85,  283.85,
  284,       284,     284,     284,
  284.45,    284.45,  284.45,  284.45,
  285,       285,     285,     285,
  285.55,    285.55,  285.55,  285.55,
  286.2,     286.2,   286.2,   286.2,
  287,       287,     287,     287,
  287.85,    287.85,  287.85,  287.85,
  288.5,     288.5,   288.5,   288.5,
  288.95,    288.95,  288.95,  288.95,
  289.5,     289.5,   289.5,   289.5,
  289.95,    289.95,  289.95,  289.95,
  290.05,    290.05,  290.05,  290.05,
  290.25,    290.25,  290.25,  290.25,
  290.05,    290.05,  290.05,  290.05,
  289.9,     289.9,   289.9,   289.9,
  290.35,    290.35,  290.35,  290.35,
  290.55,    290.55,  290.55,  290.55,
  290.4,     290.4,   290.4,   290.4,
  290.35,    290.35,  290.35,  290.35,
  290.25,    290.25,  290.25,  290.25,
  289.75,    289.75,  289.75,  289.75,
  289.2,     289.2,   289.2,   289.2,
  288.9,     288.9,   288.9,   288.9,
  289,       289,     289,     289,
  289,       289,     289,     289,
  288.65,    288.65,  288.65,  288.65,
  288.05,    288.05,  288.05,  288.05,
  287.25,    287.25,  287.25,  287.25,
  286.8,     286.8,   286.8,   286.8,
  286.45,    286.45,  286.45,  286.45,
  286.1,     286.1,   286.1,   286.1,
  286.2,     286.2,   286.2,   286.2,
  286.4,     286.4,   286.4,   286.4,
  286.3,     286.3,   286.3,   286.3,
  286.55,    286.55,  286.55,  286.55,
  287.1,     287.1,   287.1,   287.1,
  287.25,    287.25,  287.25,  287.25,
  287.45,    287.45,  287.45,  287.45,
  287.3,     287.3,   287.3,   287.3,
  286.7,     286.7,   286.7,   286.7,
  286.5,     286.5,   286.5,   286.5,
  286.55,    286.55,  286.55,  286.55,
  286.45,    286.45,  286.45,  286.45,
  286.4,     286.4,   286.4,   286.4,
  286.55,    286.55,  286.55,  286.55,
  286.8,     286.8,   286.8,   286.8,
  286.95,    286.95,  286.95,  286.95,
  286.95,    286.95,  286.95,  286.95,
  287.1,     287.1,   287.1,   287.1,
  287.35,    287.35,  287.35,  287.35,
  287.25,    287.25,  287.25,  287.25,
  287.25,    287.25,  287.25,  287.25,
  287.65,    287.65,  287.65,  287.65,
  288.05,    288.05,  288.05,  288.05,
  288.25,    288.25,  288.25,  288.25,
  288.9,     288.9,   288.9,   288.9,
  289.9,     289.9,   289.9,   289.9,
  290.6,     290.6,   290.6,   290.6,
  290.45,    290.45,  290.45,  290.45,
  288.8,     288.8,   288.8,   288.8,
  287.4,     287.4,   287.4,   287.4,
  288.35,    288.35,  288.35,  288.35,
  289.7,     289.7,   289.7,   289.7,
  289.05,    289.05,  289.05,  289.05,
  288.3,     288.3,   288.3,   288.3,
  288.8,     288.8,   288.8,   288.8,
  289.65,    289.65,  289.65,  289.65,
  290.1,     290.1,   290.1,   290.1,
  290.1,     290.1,   290.1,   290.1,
  290.1,     290.1,   290.1,   290.1,
  290,       290,     290,     290,
  289.5,     289.5,   289.5,   289.5,
  289.3,     289.3,   289.3,   289.3,
  289.45,    289.45,  289.45,  289.45,
  288.85,    288.85,  288.85,  288.85,
  287.45,    287.45,  287.45,  287.45,
  286.3,     286.3,   286.3,   286.3,
  285.75,    285.75,  285.75,  285.75,
  285.4,     285.4,   285.4,   285.4,
  285.1,     285.1,   285.1,   285.1,
  285.1,     285.1,   285.1,   285.1,
  285.15,    285.15,  285.15,  285.15,
  285.05,    285.05,  285.05,  285.05,
  284.9,     284.9,   284.9,   284.9,
  284.7,     284.7,   284.7,   284.7,
  284.55,    284.55,  284.55,  284.55,
  284.45,    284.45,  284.45,  284.45,
  284.6,     284.6,   284.6,   284.6,
  284.85,    284.85,  284.85,  284.85,
  284.7,     284.7,   284.7,   284.7,
  284.3,     284.3,   284.3,   284.3,
  284.15,    284.15,  284.15,  284.15,
  284.1,     284.1,   284.1,   284.1,
  284.1,     284.1,   284.1,   284.1,
  284.4,     284.4,   284.4,   284.4,
  284.75,    284.75,  284.75,  284.75,
  285,       285,     285,     285,
  285.35,    285.35,  285.35,  285.35,
  286.05,    286.05,  286.05,  286.05,
  286.95,    286.95,  286.95,  286.95,
  287.45,    287.45,  287.45,  287.45,
  287.7,     287.7,   287.7,   287.7,
  288.05,    288.05,  288.05,  288.05,
  288.2,     288.2,   288.2,   288.2,
  288.15,    288.15,  288.15,  288.15,
  288.35,    288.35,  288.35,  288.35,
  288.9,     288.9,   288.9,   288.9,
  289.2,     289.2,   289.2,   289.2,
  288.15,    288.15,  288.15,  288.15,
  287.6,     287.6,   287.6,   287.6,
  288.35,    288.35,  288.35,  288.35,
  289.05,    289.05,  289.05,  289.05,
  289.6,     289.6,   289.6,   289.6,
  289.9,     289.9,   289.9,   289.9,
  288.9,     288.9,   288.9,   288.9,
  286.5,     286.5,   286.5,   286.5,
  285.9,     285.9,   285.9,   285.9,
  286.35,    286.35,  286.35,  286.35,
  286.6,     286.6,   286.6,   286.6,
  286.9,     286.9,   286.9,   286.9,
  286.6,     286.6,   286.6,   286.6,
  286.1,     286.1,   286.1,   286.1,
  285.6,     285.6,   285.6,   285.6,
  285.4,     285.4,   285.4,   285.4,
  285.2,     285.2,   285.2,   285.2,
  284.9,     284.9,   284.9,   284.9,
  284.7,     284.7,   284.7,   284.7,
  284.55,    284.55,  284.55,  284.55,
  284.35,    284.35,  284.35,  284.35,
  284.25,    284.25,  284.25,  284.25,
  284.3,     284.3,   284.3,   284.3,
  284.4,     284.4,   284.4,   284.4,
  284.5,     284.5,   284.5,   284.5,
  284.5,     284.5,   284.5,   284.5,
  284.4,     284.4,   284.4,   284.4,
  284.25,    284.25,  284.25,  284.25,
  284.25,    284.25,  284.25,  284.25,
  284.25,    284.25,  284.25,  284.25,
  284.1,     284.1,   284.1,   284.1,
  284.15,    284.15,  284.15,  284.15,
  284.35,    284.35,  284.35,  284.35,
  284.55,    284.55,  284.55,  284.55,
  284.8,     284.8,   284.8,   284.8,
  285.1,     285.1,   285.1,   285.1,
  285.45,    285.45,  285.45,  285.45,
  285.85,    285.85,  285.85,  285.85,
  286.2,     286.2,   286.2,   286.2,
  286.5,     286.5,   286.5,   286.5,
  286.4,     286.4,   286.4,   286.4,
  285.9,     285.9,   285.9,   285.9,
  285.5,     285.5,   285.5,   285.5,
  285.4,     285.4,   285.4,   285.4,
  285.55,    285.55,  285.55,  285.55,
  285.65,    285.65,  285.65,  285.65,
  285.7,     285.7,   285.7,   285.7,
  285.7,     285.7,   285.7,   285.7,
  285.6,     285.6,   285.6,   285.6,
  285.6,     285.6,   285.6,   285.6,
  285.75,    285.75,  285.75,  285.75,
  285.75,    285.75,  285.75,  285.75,
  285.65,    285.65,  285.65,  285.65,
  285.65,    285.65,  285.65,  285.65,
  285.75,    285.75,  285.75,  285.75,
  285.8,     285.8,   285.8,   285.8,
  285.75,    285.75,  285.75,  285.75,
  285.85,    285.85,  285.85,  285.85,
  285.65,    285.65,  285.65,  285.65,
  285.2,     285.2,   285.2,   285.2,
  285.05,    285.05,  285.05,  285.05,
  284.95,    284.95,  284.95,  284.95,
  284.7,     284.7,   284.7,   284.7,
  284.5,     284.5,   284.5,   284.5,
  284.4,     284.4,   284.4,   284.4,
  284.35,    284.35,  284.35,  284.35,
  284.35,    284.35,  284.35,  284.35,
  284.35,    284.35,  284.35,  284.35,
  284.3,     284.3,   284.3,   284.3,
  284.25,    284.25,  284.25,  284.25,
  284.2,     284.2,   284.2,   284.2,
  284.1,     284.1,   284.1,   284.1,
  284.05,    284.05,  284.05,  284.05,
  284.05,    284.05,  284.05,  284.05,
  284.05,    284.05,  284.05,  284.05,
  284,       284,     284,     284,
  283.95,    283.95,  283.95,  283.95,
  283.95,    283.95,  283.95,  283.95,
  283.9,     283.9,   283.9,   283.9,
  283.8,     283.8,   283.8,   283.8,
  283.85,    283.85,  283.85,  283.85,
  284.05,    284.05,  284.05,  284.05,
  284.2,     284.2,   284.2,   284.2,
  284.2,     284.2,   284.2,   284.2,
  284.4,     284.4,   284.4,   284.4,
  284.85,    284.85,  284.85,  284.85,
  285.2,     285.2,   285.2,   285.2,
  285.55,    285.55,  285.55,  285.55,
  285.95,    285.95,  285.95,  285.95,
  286.2,     286.2,   286.2,   286.2,
  286.4,     286.4,   286.4,   286.4,
  286.65,    286.65,  286.65,  286.65,
  286.6,     286.6,   286.6,   286.6,
  286.55,    286.55,  286.55,  286.55,
  286.55,    286.55,  286.55,  286.55,
  286.5,     286.5,   286.5,   286.5,
  286.5,     286.5,   286.5,   286.5,
  286.6,     286.6,   286.6,   286.6,
  286.75,    286.75,  286.75,  286.75,
  286.5,     286.5,   286.5,   286.5,
  286.4,     286.4,   286.4,   286.4,
  286.7,     286.7,   286.7,   286.7,
  286.7,     286.7,   286.7,   286.7,
  286.6,     286.6,   286.6,   286.6,
  286.6,     286.6,   286.6,   286.6,
  286.4,     286.4,   286.4,   286.4,
  286.1,     286.1,   286.1,   286.1,
  285.75,    285.75,  285.75,  285.75,
  285.5,     285.5,   285.5,   285.5,
  285.35,    285.35,  285.35,  285.35,
  285.15,    285.15,  285.15,  285.15,
  284.8,     284.8,   284.8,   284.8,
  284.25,    284.25,  284.25,  284.25,
  283.75,    283.75,  283.75,  283.75,
  283.5,     283.5,   283.5,   283.5,
  283.45,    283.45,  283.45,  283.45,
  282.8,     282.8,   282.8,   282.8,
  281.85,    281.85,  281.85,  281.85,
  281.45,    281.45,  281.45,  281.45,
  281.25,    281.25,  281.25,  281.25,
  281,       281,     281,     281,
  280.6,     280.6,   280.6,   280.6,
  280.4,     280.4,   280.4,   280.4,
  280.25,    280.25,  280.25,  280.25,
  279.8,     279.8,   279.8,   279.8,
  279.1,     279.1,   279.1,   279.1,
  278.6,     278.6,   278.6,   278.6,
  278.75,    278.75,  278.75,  278.75,
  279,       279,     279,     279,
  279.25,    279.25,  279.25,  279.25,
  279.95,    279.95,  279.95,  279.95,
  281.05,    281.05,  281.05,  281.05,
  282.65,    282.65,  282.65,  282.65,
  284.25,    284.25,  284.25,  284.25,
  285.35,    285.35,  285.35,  285.35,
  286.2,     286.2,   286.2,   286.2,
  286.95,    286.95,  286.95,  286.95,
  287.6,     287.6,   287.6,   287.6,
  288.2,     288.2,   288.2,   288.2,
  288.7,     288.7,   288.7,   288.7,
  288.95,    288.95,  288.95,  288.95,
  289.25,    289.25,  289.25,  289.25,
  289.5,     289.5,   289.5,   289.5,
  289.65,    289.65,  289.65,  289.65,
  289.8,     289.8,   289.8,   289.8,
  289.85,    289.85,  289.85,  289.85,
  289.7,     289.7,   289.7,   289.7,
  289.4,     289.4,   289.4,   289.4,
  289.2,     289.2,   289.2,   289.2,
  289.05,    289.05,  289.05,  289.05,
  289.05,    289.05,  289.05,  289.05,
  289,       289,     289,     289,
  288.1,     288.1,   288.1,   288.1,
  287,       287,     287,     287,
  286.35,    286.35,  286.35,  286.35,
  285.9,     285.9,   285.9,   285.9,
  285.6,     285.6,   285.6,   285.6,
  285.35,    285.35,  285.35,  285.35,
  285.15,    285.15,  285.15,  285.15,
  285,       285,     285,     285,
  284.8,     284.8,   284.8,   284.8,
  284.55,    284.55,  284.55,  284.55,
  284.35,    284.35,  284.35,  284.35,
  284.2,     284.2,   284.2,   284.2,
  284.2,     284.2,   284.2,   284.2,
  284.25,    284.25,  284.25,  284.25,
  284.3,     284.3,   284.3,   284.3,
  284.45,    284.45,  284.45,  284.45,
  284.55,    284.55,  284.55,  284.55,
  284.55,    284.55,  284.55,  284.55,
  284.55,    284.55,  284.55,  284.55,
  284.55,    284.55,  284.55,  284.55,
  284.6,     284.6,   284.6,   284.6,
  284.7,     284.7,   284.7,   284.7,
  284.75,    284.75,  284.75,  284.75,
  284.75,    284.75,  284.75,  284.75,
  284.75,    284.75,  284.75,  284.75,
  284.8,     284.8,   284.8,   284.8,
  284.85,    284.85,  284.85,  284.85,
  284.9,     284.9,   284.9,   284.9,
  285,       285,     285,     285,
  285.2,     285.2,   285.2,   285.2,
  285.4,     285.4,   285.4,   285.4,
  285.45,    285.45,  285.45,  285.45,
  285.45,    285.45,  285.45,  285.45,
  285.55,    285.55,  285.55,  285.55,
  285.7,     285.7,   285.7,   285.7,
  285.9,     285.9,   285.9,   285.9,
  286.2,     286.2,   286.2,   286.2,
  286.6,     286.6,   286.6,   286.6,
  287.05,    287.05,  287.05,  287.05,
  287.75,    287.75,  287.75,  287.75,
  288.25,    288.25,  288.25,  288.25,
  288,       288,     288,     288,
  287.55,    287.55,  287.55,  287.55,
  287.4,     287.4,   287.4,   287.4,
  287.45,    287.45,  287.45,  287.45,
  287.55,    287.55,  287.55,  287.55,
  287.75,    287.75,  287.75,  287.75,
  287.95,    287.95,  287.95,  287.95,
  288.25,    288.25,  288.25,  288.25,
  288.75,    288.75,  288.75,  288.75,
  289.25,    289.25,  289.25,  289.25,
  289.2,     289.2,   289.2,   289.2,
  288.7,     288.7,   288.7,   288.7,
  288.25,    288.25,  288.25,  288.25,
  288.05,    288.05,  288.05,  288.05,
  287.9,     287.9,   287.9,   287.9,
  287.5,     287.5,   287.5,   287.5,
  287.15,    287.15,  287.15,  287.15,
  286.9,     286.9,   286.9,   286.9,
  286.65,    286.65,  286.65,  286.65,
  286.5,     286.5,   286.5,   286.5,
  286.3,     286.3,   286.3,   286.3,
  286.05,    286.05,  286.05,  286.05,
  285.95,    285.95,  285.95,  285.95,
  286,       286,     286,     286,
  286.1,     286.1,   286.1,   286.1,
  286.15,    286.15,  286.15,  286.15,
  286.15,    286.15,  286.15,  286.15,
  286.2,     286.2,   286.2,   286.2,
  286.25,    286.25,  286.25,  286.25,
  286.3,     286.3,   286.3,   286.3,
  286.4,     286.4,   286.4,   286.4,
  286.4,     286.4,   286.4,   286.4,
  286.4,     286.4,   286.4,   286.4,
  286.55,    286.55,  286.55,  286.55,
  286.8,     286.8,   286.8,   286.8,
  287.05,    287.05,  287.05,  287.05,
  287.25,    287.25,  287.25,  287.25,
  287.45,    287.45,  287.45,  287.45,
  287.7,     287.7,   287.7,   287.7,
  288,       288,     288,     288,
  288.4,     288.4,   288.4,   288.4,
  289.1,     289.1,   289.1,   289.1,
  289.9,     289.9,   289.9,   289.9,
  290.55,    290.55,  290.55,  290.55,
  291.35,    291.35,  291.35,  291.35,
  292.05,    292.05,  292.05,  292.05,
  292.35,    292.35,  292.35,  292.35,
  292.45,    292.45,  292.45,  292.45,
  292.35,    292.35,  292.35,  292.35,
  291.55,    291.55,  291.55,  291.55,
  288.65,    288.65,  288.65,  288.65,
  285.95,    285.95,  285.95,  285.95,
  285.25,    285.25,  285.25,  285.25,
  285.25,    285.25,  285.25,  285.25,
  285.6,     285.6,   285.6,   285.6,
  285.9,     285.9,   285.9,   285.9,
  286.3,     286.3,   286.3,   286.3,
  286.95,    286.95,  286.95,  286.95,
  287.5,     287.5,   287.5,   287.5,
  287.7,     287.7,   287.7,   287.7,
  287.45,    287.45,  287.45,  287.45,
  286.8,     286.8,   286.8,   286.8,
  286,       286,     286,     286,
  285.25,    285.25,  285.25,  285.25,
  284.8,     284.8,   284.8,   284.8,
  284.45,    284.45,  284.45,  284.45,
  284.15,    284.15,  284.15,  284.15,
  284,       284,     284,     284,
  283.95,    283.95,  283.95,  283.95,
  283.95,    283.95,  283.95,  283.95,
  283.9,     283.9,   283.9,   283.9,
  283.65,    283.65,  283.65,  283.65,
  283.3,     283.3,   283.3,   283.3,
  283.4,     283.4,   283.4,   283.4,
  283.85,    283.85,  283.85,  283.85,
  284.15,    284.15,  284.15,  284.15,
  284.2,     284.2,   284.2,   284.2,
  284.1,     284.1,   284.1,   284.1,
  284.05,    284.05,  284.05,  284.05,
  284.2,     284.2,   284.2,   284.2,
  284.65,    284.65,  284.65,  284.65,
  285.1,     285.1,   285.1,   285.1,
  285.6,     285.6,   285.6,   285.6,
  286.3,     286.3,   286.3,   286.3,
  287,       287,     287,     287,
  287.3,     287.3,   287.3,   287.3,
  287.5,     287.5,   287.5,   287.5,
  288.05,    288.05,  288.05,  288.05,
  288.35,    288.35,  288.35,  288.35,
  288.65,    288.65,  288.65,  288.65,
  288.7,     288.7,   288.7,   288.7,
  289.2,     289.2,   289.2,   289.2,
  290.2,     290.2,   290.2,   290.2,
  290.3,     290.3,   290.3,   290.3,
  289.35,    289.35,  289.35,  289.35,
  289,       289,     289,     289,
  289.15,    289.15,  289.15,  289.15,
  289.4,     289.4,   289.4,   289.4,
  289.85,    289.85,  289.85,  289.85,
  290.05,    290.05,  290.05,  290.05,
  290.4,     290.4,   290.4,   290.4,
  290.25,    290.25,  290.25,  290.25,
  290.85,    290.85,  290.85,  290.85,
  291.55,    291.55,  291.55,  291.55,
  291.45,    291.45,  291.45,  291.45,
  291.7,     291.7,   291.7,   291.7,
  292.25,    292.25,  292.25,  292.25,
  292.4,     292.4,   292.4,   292.4,
  292.05,    292.05,  292.05,  292.05,
  291.7,     291.7,   291.7,   291.7,
  291.25,    291.25,  291.25,  291.25,
  290.55,    290.55,  290.55,  290.55,
  289.65,    289.65,  289.65,  289.65,
  288.8,     288.8,   288.8,   288.8,
  288.3,     288.3,   288.3,   288.3,
  287.9,     287.9,   287.9,   287.9,
  287.3,     287.3,   287.3,   287.3,
  286.6,     286.6,   286.6,   286.6,
  286.1,     286.1,   286.1,   286.1,
  285.55,    285.55,  285.55,  285.55,
  285.35,    285.35,  285.35,  285.35,
  285.2,     285.2,   285.2,   285.2,
  284.95,    284.95,  284.95,  284.95,
  285.1,     285.1,   285.1,   285.1,
  285.3,     285.3,   285.3,   285.3,
  285.4,     285.4,   285.4,   285.4,
  285.35,    285.35,  285.35,  285.35,
  285.45,    285.45,  285.45,  285.45,
  286.05,    286.05,  286.05,  286.05,
  287.15,    287.15,  287.15,  287.15,
  287.95,    287.95,  287.95,  287.95,
  288.35,    288.35,  288.35,  288.35,
  288.9,     288.9,   288.9,   288.9,
  289.65,    289.65,  289.65,  289.65,
  290.45,    290.45,  290.45,  290.45,
  291.3,     291.3,   291.3,   291.3,
  292.4,     292.4,   292.4,   292.4,
  293.5,     293.5,   293.5,   293.5,
  294.3,     294.3,   294.3,   294.3,
  294.9,     294.9,   294.9,   294.9,
  295.3,     295.3,   295.3,   295.3,
  295.25,    295.25,  295.25,  295.25,
  294.45,    294.45,  294.45,  294.45,
  292.2,     292.2,   292.2,   292.2,
  290,       290,     290,     290,
  289.3,     289.3,   289.3,   289.3,
  289.05,    289.05,  289.05,  289.05,
  289.05,    289.05,  289.05,  289.05,
  289.3,     289.3,   289.3,   289.3,
  289.3,     289.3,   289.3,   289.3,
  289.15,    289.15,  289.15,  289.15,
  289.15,    289.15,  289.15,  289.15,
  289.15,    289.15,  289.15,  289.15,
  289.2,     289.2,   289.2,   289.2,
  289.3,     289.3,   289.3,   289.3,
  289.3,     289.3,   289.3,   289.3,
  288.85,    288.85,  288.85,  288.85,
  288.4,     288.4,   288.4,   288.4,
  288.35,    288.35,  288.35,  288.35,
  288.3,     288.3,   288.3,   288.3,
  288.2,     288.2,   288.2,   288.2,
  288.15,    288.15,  288.15,  288.15,
  288.15,    288.15,  288.15,  288.15,
  288.15,    288.15,  288.15,  288.15,
  288.15,    288.15,  288.15,  288.15,
  288.15,    288.15,  288.15,  288.15,
  288.15,    288.15,  288.15,  288.15,
  288.1,     288.1,   288.1,   288.1,
  287.95,    287.95,  287.95,  287.95,
  287.75,    287.75,  287.75,  287.75,
  287.55,    287.55,  287.55,  287.55,
  287.45,    287.45,  287.45,  287.45,
  287.45,    287.45,  287.45,  287.45,
  287.4,     287.4,   287.4,   287.4,
  287.35,    287.35,  287.35,  287.35,
  287.25,    287.25,  287.25,  287.25,
  287.1,     287.1,   287.1,   287.1,
  287.1,     287.1,   287.1,   287.1,
  287.2,     287.2,   287.2,   287.2,
  287.3,     287.3,   287.3,   287.3,
  287.45,    287.45,  287.45,  287.45,
  287.55,    287.55,  287.55,  287.55,
  287.55,    287.55,  287.55,  287.55,
  287.6,     287.6,   287.6,   287.6,
  287.75,    287.75,  287.75,  287.75,
  288,       288,     288,     288,
  288.1,     288.1,   288.1,   288.1,
  288,       288,     288,     288,
  288,       288,     288,     288,
  288.05,    288.05,  288.05,  288.05,
  288.1,     288.1,   288.1,   288.1,
  288.2,     288.2,   288.2,   288.2,
  288.35,    288.35,  288.35,  288.35,
  288.3,     288.3,   288.3,   288.3,
  288.15,    288.15,  288.15,  288.15,
  288.15,    288.15,  288.15,  288.15,
  288.2,     288.2,   288.2,   288.2,
  288.25,    288.25,  288.25,  288.25,
  288.05,    288.05,  288.05,  288.05,
  287.75,    287.75,  287.75,  287.75,
  287.35,    287.35,  287.35,  287.35,
  286.9,     286.9,   286.9,   286.9,
  286.5,     286.5,   286.5,   286.5,
  285.9,     285.9,   285.9,   285.9,
  285.55,    285.55,  285.55,  285.55,
  285.6,     285.6,   285.6,   285.6,
  285.6,     285.6,   285.6,   285.6,
  285.55,    285.55,  285.55,  285.55,
  285.55,    285.55,  285.55,  285.55,
  285.5,     285.5,   285.5,   285.5,
  285.45,    285.45,  285.45,  285.45,
  285.45,    285.45,  285.45,  285.45,
  285.45,    285.45,  285.45,  285.45,
  285.45,    285.45,  285.45,  285.45,
  285.45,    285.45,  285.45,  285.45,
  285.4,     285.4,   285.4,   285.4,
  285.25,    285.25,  285.25,  285.25,
  284.85,    284.85,  284.85,  284.85,
  284.4,     284.4,   284.4,   284.4,
  284.1,     284.1,   284.1,   284.1,
  283.9,     283.9,   283.9,   283.9,
  283.8,     283.8,   283.8,   283.8,
  283.75,    283.75,  283.75,  283.75,
  283.8,     283.8,   283.8,   283.8,
  284.15,    284.15,  284.15,  284.15,
  284.65,    284.65,  284.65,  284.65,
  284.9,     284.9,   284.9,   284.9,
  285.15,    285.15,  285.15,  285.15,
  285.55,    285.55,  285.55,  285.55,
  285.9,     285.9,   285.9,   285.9,
  286.4,     286.4,   286.4,   286.4,
  287.05,    287.05,  287.05,  287.05,
  287.5,     287.5,   287.5,   287.5,
  287.7,     287.7,   287.7,   287.7,
  287.9,     287.9,   287.9,   287.9,
  288.15,    288.15,  288.15,  288.15,
  288.45,    288.45,  288.45,  288.45,
  289.05,    289.05,  289.05,  289.05,
  289.7,     289.7,   289.7,   289.7,
  290.1,     290.1,   290.1,   290.1,
  290.6,     290.6,   290.6,   290.6,
  291.45,    291.45,  291.45,  291.45,
  291.95,    291.95,  291.95,  291.95,
  292.15,    292.15,  292.15,  292.15,
  292.3,     292.3,   292.3,   292.3,
  292.25,    292.25,  292.25,  292.25,
  290.35,    290.35,  290.35,  290.35,
  287.55,    287.55,  287.55,  287.55,
  287.15,    287.15,  287.15,  287.15,
  288.05,    288.05,  288.05,  288.05,
  288.75,    288.75,  288.75,  288.75,
  288.8,     288.8,   288.8,   288.8,
  288.35,    288.35,  288.35,  288.35,
  287.85,    287.85,  287.85,  287.85,
  287.4,     287.4,   287.4,   287.4,
  287.25,    287.25,  287.25,  287.25,
  287,       287,     287,     287,
  286.5,     286.5,   286.5,   286.5,
  286.05,    286.05,  286.05,  286.05,
  285.7,     285.7,   285.7,   285.7,
  285.3,     285.3,   285.3,   285.3,
  285.15,    285.15,  285.15,  285.15,
  285.1,     285.1,   285.1,   285.1,
  284.85,    284.85,  284.85,  284.85,
  284.25,    284.25,  284.25,  284.25,
  283.4,     283.4,   283.4,   283.4,
  282.95,    282.95,  282.95,  282.95,
  282.75,    282.75,  282.75,  282.75,
  282.55,    282.55,  282.55,  282.55,
  282.45,    282.45,  282.45,  282.45,
  282.3,     282.3,   282.3,   282.3,
  282.3,     282.3,   282.3,   282.3,
  282.75,    282.75,  282.75,  282.75,
  283.3,     283.3,   283.3,   283.3,
  284,       284,     284,     284,
  284.95,    284.95,  284.95,  284.95,
  286.1,     286.1,   286.1,   286.1,
  287.2,     287.2,   287.2,   287.2,
  288.05,    288.05,  288.05,  288.05,
  288.6,     288.6,   288.6,   288.6,
  289,       289,     289,     289,
  289.7,     289.7,   289.7,   289.7,
  290.55,    290.55,  290.55,  290.55,
  291.15,    291.15,  291.15,  291.15,
  291.55,    291.55,  291.55,  291.55,
  292,       292,     292,     292,
  292.55,    292.55,  292.55,  292.55,
  293,       293,     293,     293,
  293.15,    293.15,  293.15,  293.15,
  292.95,    292.95,  292.95,  292.95,
  292.7,     292.7,   292.7,   292.7,
  292.5,     292.5,   292.5,   292.5,
  292.25,    292.25,  292.25,  292.25,
  292.1,     292.1,   292.1,   292.1,
  291.7,     291.7,   291.7,   291.7,
  290.55,    290.55,  290.55,  290.55,
  289.3,     289.3,   289.3,   289.3,
  288.65,    288.65,  288.65,  288.65,
  288.4,     288.4,   288.4,   288.4,
  288.45,    288.45,  288.45,  288.45,
  288.55,    288.55,  288.55,  288.55,
  288.45,    288.45,  288.45,  288.45,
  288.3,     288.3,   288.3,   288.3,
  288.3,     288.3,   288.3,   288.3,
  288.45,    288.45,  288.45,  288.45,
  288.6,     288.6,   288.6,   288.6,
  288.35,    288.35,  288.35,  288.35,
  287.55,    287.55,  287.55,  287.55,
  286.85,    286.85,  286.85,  286.85,
  286.45,    286.45,  286.45,  286.45,
  286.1,     286.1,   286.1,   286.1,
  285.85,    285.85,  285.85,  285.85,
  285.55,    285.55,  285.55,  285.55,
  285.05,    285.05,  285.05,  285.05,
  284.5,     284.5,   284.5,   284.5,
  284.15,    284.15,  284.15,  284.15,
  283.9,     283.9,   283.9,   283.9,
  283.65,    283.65,  283.65,  283.65,
  283.5,     283.5,   283.5,   283.5,
  283.5,     283.5,   283.5,   283.5,
  283.85,    283.85,  283.85,  283.85,
  284.6,     284.6,   284.6,   284.6,
  285.4,     285.4,   285.4,   285.4,
  286.05,    286.05,  286.05,  286.05,
  286.7,     286.7,   286.7,   286.7,
  287.35,    287.35,  287.35,  287.35,
  288.05,    288.05,  288.05,  288.05,
  288.8,     288.8,   288.8,   288.8,
  289.4,     289.4,   289.4,   289.4,
  289.65,    289.65,  289.65,  289.65,
  290.1,     290.1,   290.1,   290.1,
  290.55,    290.55,  290.55,  290.55,
  290.6,     290.6,   290.6,   290.6,
  290.9,     290.9,   290.9,   290.9,
  291.25,    291.25,  291.25,  291.25,
  291.5,     291.5,   291.5,   291.5,
  291.55,    291.55,  291.55,  291.55,
  291.3,     291.3,   291.3,   291.3,
  291.35,    291.35,  291.35,  291.35,
  291.65,    291.65,  291.65,  291.65,
  291.75,    291.75,  291.75,  291.75,
  291.7,     291.7,   291.7,   291.7,
  291.75,    291.75,  291.75,  291.75,
  291.75,    291.75,  291.75,  291.75,
  291.6,     291.6,   291.6,   291.6,
  291.55,    291.55,  291.55,  291.55,
  291.25,    291.25,  291.25,  291.25,
  289.8,     289.8,   289.8,   289.8,
  288,       288,     288,     288,
  287.35,    287.35,  287.35,  287.35,
  287.3,     287.3,   287.3,   287.3,
  286.95,    286.95,  286.95,  286.95,
  286.4,     286.4,   286.4,   286.4,
  286.05,    286.05,  286.05,  286.05,
  285.95,    285.95,  285.95,  285.95,
  285.85,    285.85,  285.85,  285.85,
  285.7,     285.7,   285.7,   285.7,
  285.6,     285.6,   285.6,   285.6,
  285.45,    285.45,  285.45,  285.45,
  285.1,     285.1,   285.1,   285.1,
  284.8,     284.8,   284.8,   284.8,
  284.5,     284.5,   284.5,   284.5,
  284.15,    284.15,  284.15,  284.15,
  283.95,    283.95,  283.95,  283.95,
  283.65,    283.65,  283.65,  283.65,
  283.3,     283.3,   283.3,   283.3,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  283.35,    283.35,  283.35,  283.35,
  283.9,     283.9,   283.9,   283.9,
  285,       285,     285,     285,
  286.35,    286.35,  286.35,  286.35,
  287.25,    287.25,  287.25,  287.25,
  287.85,    287.85,  287.85,  287.85,
  288.45,    288.45,  288.45,  288.45,
  289.15,    289.15,  289.15,  289.15,
  290,       290,     290,     290,
  290.7,     290.7,   290.7,   290.7,
  291.1,     291.1,   291.1,   291.1,
  291.5,     291.5,   291.5,   291.5,
  291.7,     291.7,   291.7,   291.7,
  291.8,     291.8,   291.8,   291.8,
  291.6,     291.6,   291.6,   291.6,
  290.15,    290.15,  290.15,  290.15,
  290.25,    290.25,  290.25,  290.25,
  292,       292,     292,     292,
  292.8,     292.8,   292.8,   292.8,
  293.15,    293.15,  293.15,  293.15,
  293.35,    293.35,  293.35,  293.35,
  293.4,     293.4,   293.4,   293.4,
  293.5,     293.5,   293.5,   293.5,
  293.3,     293.3,   293.3,   293.3,
  292.7,     292.7,   292.7,   292.7,
  291.55,    291.55,  291.55,  291.55,
  290.3,     290.3,   290.3,   290.3,
  289.8,     289.8,   289.8,   289.8,
  289.45,    289.45,  289.45,  289.45,
  289.1,     289.1,   289.1,   289.1,
  288.8,     288.8,   288.8,   288.8,
  288.45,    288.45,  288.45,  288.45,
  288.05,    288.05,  288.05,  288.05,
  287.85,    287.85,  287.85,  287.85,
  287.85,    287.85,  287.85,  287.85,
  287.65,    287.65,  287.65,  287.65,
  287.1,     287.1,   287.1,   287.1,
  286.9,     286.9,   286.9,   286.9,
  287,       287,     287,     287,
  286.85,    286.85,  286.85,  286.85,
  286.5,     286.5,   286.5,   286.5,
  286.35,    286.35,  286.35,  286.35,
  286.4,     286.4,   286.4,   286.4,
  286.15,    286.15,  286.15,  286.15,
  285.95,    285.95,  285.95,  285.95,
  285.9,     285.9,   285.9,   285.9,
  286,       286,     286,     286,
  286.1,     286.1,   286.1,   286.1,
  286,       286,     286,     286,
  286.3,     286.3,   286.3,   286.3,
  287.05,    287.05,  287.05,  287.05,
  287.65,    287.65,  287.65,  287.65,
  288.1,     288.1,   288.1,   288.1,
  288.75,    288.75,  288.75,  288.75,
  289.45,    289.45,  289.45,  289.45,
  290,       290,     290,     290,
  290.6,     290.6,   290.6,   290.6,
  291.5,     291.5,   291.5,   291.5,
  291.9,     291.9,   291.9,   291.9,
  291.7,     291.7,   291.7,   291.7,
  291.95,    291.95,  291.95,  291.95,
  292,       292,     292,     292,
  290.65,    290.65,  290.65,  290.65,
  289.1,     289.1,   289.1,   289.1,
  288.55,    288.55,  288.55,  288.55,
  288.75,    288.75,  288.75,  288.75,
  289.05,    289.05,  289.05,  289.05,
  288.65,    288.65,  288.65,  288.65,
  288.15,    288.15,  288.15,  288.15,
  288.2,     288.2,   288.2,   288.2,
  288.8,     288.8,   288.8,   288.8,
  289.75,    289.75,  289.75,  289.75,
  290.1,     290.1,   290.1,   290.1,
  290,       290,     290,     290,
  290.05,    290.05,  290.05,  290.05,
  289.75,    289.75,  289.75,  289.75,
  289.3,     289.3,   289.3,   289.3,
  288.95,    288.95,  288.95,  288.95,
  288.35,    288.35,  288.35,  288.35,
  287.6,     287.6,   287.6,   287.6,
  286.85,    286.85,  286.85,  286.85,
  286.3,     286.3,   286.3,   286.3,
  286.05,    286.05,  286.05,  286.05,
  285.8,     285.8,   285.8,   285.8,
  285.25,    285.25,  285.25,  285.25,
  284.8,     284.8,   284.8,   284.8,
  284.9,     284.9,   284.9,   284.9,
  285,       285,     285,     285,
  284.75,    284.75,  284.75,  284.75,
  284.4,     284.4,   284.4,   284.4,
  284.1,     284.1,   284.1,   284.1,
  283.75,    283.75,  283.75,  283.75,
  283.45,    283.45,  283.45,  283.45,
  283.4,     283.4,   283.4,   283.4,
  283.55,    283.55,  283.55,  283.55,
  283.75,    283.75,  283.75,  283.75,
  283.95,    283.95,  283.95,  283.95,
  284.15,    284.15,  284.15,  284.15,
  284.55,    284.55,  284.55,  284.55,
  285.45,    285.45,  285.45,  285.45,
  286.65,    286.65,  286.65,  286.65,
  287.55,    287.55,  287.55,  287.55,
  287.9,     287.9,   287.9,   287.9,
  288.25,    288.25,  288.25,  288.25,
  288.7,     288.7,   288.7,   288.7,
  288.75,    288.75,  288.75,  288.75,
  288.7,     288.7,   288.7,   288.7,
  288.75,    288.75,  288.75,  288.75,
  288.55,    288.55,  288.55,  288.55,
  288.65,    288.65,  288.65,  288.65,
  288.9,     288.9,   288.9,   288.9,
  288.65,    288.65,  288.65,  288.65,
  288.35,    288.35,  288.35,  288.35,
  288.1,     288.1,   288.1,   288.1,
  287.8,     287.8,   287.8,   287.8,
  287.45,    287.45,  287.45,  287.45,
  287.15,    287.15,  287.15,  287.15,
  287.1,     287.1,   287.1,   287.1,
  287.3,     287.3,   287.3,   287.3,
  287.6,     287.6,   287.6,   287.6,
  288,       288,     288,     288,
  288.25,    288.25,  288.25,  288.25,
  288.35,    288.35,  288.35,  288.35,
  288.6,     288.6,   288.6,   288.6,
  288.85,    288.85,  288.85,  288.85,
  289,       289,     289,     289,
  289.05,    289.05,  289.05,  289.05,
  288.75,    288.75,  288.75,  288.75,
  288.2,     288.2,   288.2,   288.2,
  288,       288,     288,     288,
  288.1,     288.1,   288.1,   288.1,
  288.1,     288.1,   288.1,   288.1,
  288,       288,     288,     288,
  287.95,    287.95,  287.95,  287.95,
  287.85,    287.85,  287.85,  287.85,
  287.7,     287.7,   287.7,   287.7,
  287.55,    287.55,  287.55,  287.55,
  287.4,     287.4,   287.4,   287.4,
  287.3,     287.3,   287.3,   287.3,
  287.2,     287.2,   287.2,   287.2,
  287.1,     287.1,   287.1,   287.1,
  287.05,    287.05,  287.05,  287.05,
  286.95,    286.95,  286.95,  286.95,
  286.8,     286.8,   286.8,   286.8,
  286.8,     286.8,   286.8,   286.8,
  286.85,    286.85,  286.85,  286.85,
  286.85,    286.85,  286.85,  286.85,
  286.85,    286.85,  286.85,  286.85,
  286.85,    286.85,  286.85,  286.85,
  287.3,     287.3,   287.3,   287.3,
  288.35,    288.35,  288.35,  288.35,
  289.55,    289.55,  289.55,  289.55,
  290.25,    290.25,  290.25,  290.25,
  290.75,    290.75,  290.75,  290.75,
  291.45,    291.45,  291.45,  291.45,
  292.25,    292.25,  292.25,  292.25,
  292.75,    292.75,  292.75,  292.75,
  292.8,     292.8,   292.8,   292.8,
  293.1,     293.1,   293.1,   293.1,
  293.2,     293.2,   293.2,   293.2,
  293.1,     293.1,   293.1,   293.1,
  293.2,     293.2,   293.2,   293.2,
  293.45,    293.45,  293.45,  293.45,
  293.7,     293.7,   293.7,   293.7,
  293.75,    293.75,  293.75,  293.75,
  293.95,    293.95,  293.95,  293.95,
  294.05,    294.05,  294.05,  294.05,
  294,       294,     294,     294,
  293.9,     293.9,   293.9,   293.9,
  293.45,    293.45,  293.45,  293.45,
  292.95,    292.95,  292.95,  292.95,
  292.5,     292.5,   292.5,   292.5,
  292,       292,     292,     292,
  291.4,     291.4,   291.4,   291.4,
  290.7,     290.7,   290.7,   290.7,
  290,       290,     290,     290,
  289.35,    289.35,  289.35,  289.35,
  288.8,     288.8,   288.8,   288.8,
  288.3,     288.3,   288.3,   288.3,
  288,       288,     288,     288,
  287.75,    287.75,  287.75,  287.75,
  287.7,     287.7,   287.7,   287.7,
  287.85,    287.85,  287.85,  287.85,
  287.7,     287.7,   287.7,   287.7,
  287.45,    287.45,  287.45,  287.45,
  287.15,    287.15,  287.15,  287.15,
  286.85,    286.85,  286.85,  286.85,
  286.7,     286.7,   286.7,   286.7,
  286.6,     286.6,   286.6,   286.6,
  286.75,    286.75,  286.75,  286.75,
  287.15,    287.15,  287.15,  287.15,
  287.45,    287.45,  287.45,  287.45,
  287.6,     287.6,   287.6,   287.6,
  287.8,     287.8,   287.8,   287.8,
  288.15,    288.15,  288.15,  288.15,
  288.45,    288.45,  288.45,  288.45,
  288.65,    288.65,  288.65,  288.65,
  288.9,     288.9,   288.9,   288.9,
  289.05,    289.05,  289.05,  289.05,
  289.1,     289.1,   289.1,   289.1,
  289.05,    289.05,  289.05,  289.05,
  289,       289,     289,     289,
  289.15,    289.15,  289.15,  289.15,
  289.3,     289.3,   289.3,   289.3,
  289.65,    289.65,  289.65,  289.65,
  290.2,     290.2,   290.2,   290.2,
  290.7,     290.7,   290.7,   290.7,
  291.25,    291.25,  291.25,  291.25,
  291.85,    291.85,  291.85,  291.85,
  292.35,    292.35,  292.35,  292.35,
  292.8,     292.8,   292.8,   292.8,
  293.1,     293.1,   293.1,   293.1,
  293.1,     293.1,   293.1,   293.1,
  293.2,     293.2,   293.2,   293.2,
  293.4,     293.4,   293.4,   293.4,
  293.65,    293.65,  293.65,  293.65,
  293.9,     293.9,   293.9,   293.9,
  293.65,    293.65,  293.65,  293.65,
  293.3,     293.3,   293.3,   293.3,
  293.15,    293.15,  293.15,  293.15,
  292.95,    292.95,  292.95,  292.95,
  292.5,     292.5,   292.5,   292.5,
  291.65,    291.65,  291.65,  291.65,
  290.75,    290.75,  290.75,  290.75,
  290.05,    290.05,  290.05,  290.05,
  289.4,     289.4,   289.4,   289.4,
  288.8,     288.8,   288.8,   288.8,
  288.25,    288.25,  288.25,  288.25,
  287.65,    287.65,  287.65,  287.65,
  287.25,    287.25,  287.25,  287.25,
  287.25,    287.25,  287.25,  287.25,
  287.4,     287.4,   287.4,   287.4,
  287.5,     287.5,   287.5,   287.5,
  287.6,     287.6,   287.6,   287.6,
  287.65,    287.65,  287.65,  287.65,
  287.6,     287.6,   287.6,   287.6,
  287.45,    287.45,  287.45,  287.45,
  287.3,     287.3,   287.3,   287.3,
  287.25,    287.25,  287.25,  287.25,
  287.25,    287.25,  287.25,  287.25,
  287.2,     287.2,   287.2,   287.2,
  287.15,    287.15,  287.15,  287.15,
  287.25,    287.25,  287.25,  287.25,
  287.4,     287.4,   287.4,   287.4,
  287.6,     287.6,   287.6,   287.6,
  288,       288,     288,     288,
  288.45,    288.45,  288.45,  288.45,
  288.7,     288.7,   288.7,   288.7,
  289,       289,     289,     289,
  289.3,     289.3,   289.3,   289.3,
  289.4,     289.4,   289.4,   289.4,
  289.5,     289.5,   289.5,   289.5,
  289.65,    289.65,  289.65,  289.65,
  289.9,     289.9,   289.9,   289.9,
  290.4,     290.4,   290.4,   290.4,
  290.85,    290.85,  290.85,  290.85,
  291.2,     291.2,   291.2,   291.2,
  291.4,     291.4,   291.4,   291.4,
  291.45,    291.45,  291.45,  291.45,
  291.85,    291.85,  291.85,  291.85,
  292.2,     292.2,   292.2,   292.2,
  292.5,     292.5,   292.5,   292.5,
  292.75,    292.75,  292.75,  292.75,
  292.8,     292.8,   292.8,   292.8,
  292.95,    292.95,  292.95,  292.95,
  293.05,    293.05,  293.05,  293.05,
  292.8,     292.8,   292.8,   292.8,
  292.35,    292.35,  292.35,  292.35,
  291.95,    291.95,  291.95,  291.95,
  291.35,    291.35,  291.35,  291.35,
  290.5,     290.5,   290.5,   290.5,
  289.55,    289.55,  289.55,  289.55,
  288.65,    288.65,  288.65,  288.65,
  287.85,    287.85,  287.85,  287.85,
  287.15,    287.15,  287.15,  287.15,
  286.55,    286.55,  286.55,  286.55,
  286,       286,     286,     286,
  285.5,     285.5,   285.5,   285.5,
  285.15,    285.15,  285.15,  285.15,
  284.95,    284.95,  284.95,  284.95,
  284.7,     284.7,   284.7,   284.7,
  284.5,     284.5,   284.5,   284.5,
  284.35,    284.35,  284.35,  284.35,
  284.15,    284.15,  284.15,  284.15,
  284.1,     284.1,   284.1,   284.1,
  284.2,     284.2,   284.2,   284.2,
  284.2,     284.2,   284.2,   284.2,
  284.55,    284.55,  284.55,  284.55,
  285.25,    285.25,  285.25,  285.25,
  285.8,     285.8,   285.8,   285.8,
  286.15,    286.15,  286.15,  286.15,
  286.4,     286.4,   286.4,   286.4,
  286.65,    286.65,  286.65,  286.65,
  286.9,     286.9,   286.9,   286.9,
  287.25,    287.25,  287.25,  287.25,
  288.2,     288.2,   288.2,   288.2,
  289.8,     289.8,   289.8,   289.8,
  291.3,     291.3,   291.3,   291.3,
  292.25,    292.25,  292.25,  292.25,
  292.7,     292.7,   292.7,   292.7,
  293.1,     293.1,   293.1,   293.1,
  293.7,     293.7,   293.7,   293.7,
  294.3,     294.3,   294.3,   294.3,
  294.6,     294.6,   294.6,   294.6,
  294.7,     294.7,   294.7,   294.7,
  295.25,    295.25,  295.25,  295.25,
  295.55,    295.55,  295.55,  295.55,
  295.3,     295.3,   295.3,   295.3,
  295.5,     295.5,   295.5,   295.5,
  295.8,     295.8,   295.8,   295.8,
  295.8,     295.8,   295.8,   295.8,
  296,       296,     296,     296,
  296.1,     296.1,   296.1,   296.1,
  296,       296,     296,     296,
  295.6,     295.6,   295.6,   295.6,
  295.25,    295.25,  295.25,  295.25,
  295.15,    295.15,  295.15,  295.15,
  294.55,    294.55,  294.55,  294.55,
  293.8,     293.8,   293.8,   293.8,
  292.85,    292.85,  292.85,  292.85,
  291.85,    291.85,  291.85,  291.85,
  291.2,     291.2,   291.2,   291.2,
  290.7,     290.7,   290.7,   290.7,
  290.25,    290.25,  290.25,  290.25,
  290,       290,     290,     290,
  289.85,    289.85,  289.85,  289.85,
  289.5,     289.5,   289.5,   289.5,
  289,       289,     289,     289,
  288.6,     288.6,   288.6,   288.6,
  288.4,     288.4,   288.4,   288.4,
  288.3,     288.3,   288.3,   288.3,
  288.2,     288.2,   288.2,   288.2,
  288.05,    288.05,  288.05,  288.05,
  287.9,     287.9,   287.9,   287.9,
  287.8,     287.8,   287.8,   287.8,
  287.75,    287.75,  287.75,  287.75,
  288.05,    288.05,  288.05,  288.05,
  288.75,    288.75,  288.75,  288.75,
  289.6,     289.6,   289.6,   289.6,
  290.5,     290.5,   290.5,   290.5,
  291.55,    291.55,  291.55,  291.55,
  292.7,     292.7,   292.7,   292.7,
  293.9,     293.9,   293.9,   293.9,
  294.9,     294.9,   294.9,   294.9,
  295.65,    295.65,  295.65,  295.65,
  296.35,    296.35,  296.35,  296.35,
  296.75,    296.75,  296.75,  296.75,
  297,       297,     297,     297,
  297.25,    297.25,  297.25,  297.25,
  297.65,    297.65,  297.65,  297.65,
  297.85,    297.85,  297.85,  297.85,
  297.9,     297.9,   297.9,   297.9,
  298.35,    298.35,  298.35,  298.35,
  298.45,    298.45,  298.45,  298.45,
  298.4,     298.4,   298.4,   298.4,
  298.6,     298.6,   298.6,   298.6,
  298.4,     298.4,   298.4,   298.4,
  298.3,     298.3,   298.3,   298.3,
  298.6,     298.6,   298.6,   298.6,
  298.45,    298.45,  298.45,  298.45,
  298.2,     298.2,   298.2,   298.2,
  298.25,    298.25,  298.25,  298.25,
  298.2,     298.2,   298.2,   298.2,
  297.9,     297.9,   297.9,   297.9,
  297.3,     297.3,   297.3,   297.3,
  296.5,     296.5,   296.5,   296.5,
  295.6,     295.6,   295.6,   295.6,
  294.65,    294.65,  294.65,  294.65,
  293.75,    293.75,  293.75,  293.75,
  292.9,     292.9,   292.9,   292.9,
  292.35,    292.35,  292.35,  292.35,
  292.25,    292.25,  292.25,  292.25,
  292.25,    292.25,  292.25,  292.25,
  292.1,     292.1,   292.1,   292.1,
  291.75,    291.75,  291.75,  291.75,
  291.35,    291.35,  291.35,  291.35,
  291.05,    291.05,  291.05,  291.05,
  290.85,    290.85,  290.85,  290.85,
  290.65,    290.65,  290.65,  290.65,
  290.6,     290.6,   290.6,   290.6,
  290.65,    290.65,  290.65,  290.65,
  290.7,     290.7,   290.7,   290.7,
  290.8,     290.8,   290.8,   290.8,
  290.55,    290.55,  290.55,  290.55,
  290.1,     290.1,   290.1,   290.1,
  290.05,    290.05,  290.05,  290.05,
  290.25,    290.25,  290.25,  290.25,
  290.5,     290.5,   290.5,   290.5,
  290.9,     290.9,   290.9,   290.9,
  291.7,     291.7,   291.7,   291.7,
  293.05,    293.05,  293.05,  293.05,
  294.15,    294.15,  294.15,  294.15,
  295.1,     295.1,   295.1,   295.1,
  296.7,     296.7,   296.7,   296.7,
  298,       298,     298,     298,
  298.2,     298.2,   298.2,   298.2,
  298.35,    298.35,  298.35,  298.35,
  298.75,    298.75,  298.75,  298.75,
  299.05,    299.05,  299.05,  299.05,
  299.25,    299.25,  299.25,  299.25,
  299.4,     299.4,   299.4,   299.4,
  299.2,     299.2,   299.2,   299.2,
  298.6,     298.6,   298.6,   298.6,
  298.4,     298.4,   298.4,   298.4,
  298.45,    298.45,  298.45,  298.45,
  298.15,    298.15,  298.15,  298.15,
  297.85,    297.85,  297.85,  297.85,
  297.85,    297.85,  297.85,  297.85,
  297.85,    297.85,  297.85,  297.85,
  297.6,     297.6,   297.6,   297.6,
  297.05,    297.05,  297.05,  297.05,
  296.35,    296.35,  296.35,  296.35,
  295.55,    295.55,  295.55,  295.55,
  294.6,     294.6,   294.6,   294.6,
  293.6,     293.6,   293.6,   293.6,
  292.65,    292.65,  292.65,  292.65,
  291.9,     291.9,   291.9,   291.9,
  291.45,    291.45,  291.45,  291.45,
  291.15,    291.15,  291.15,  291.15,
  290.9,     290.9,   290.9,   290.9,
  290.7,     290.7,   290.7,   290.7,
  290.45,    290.45,  290.45,  290.45,
  290.05,    290.05,  290.05,  290.05,
  289.75,    289.75,  289.75,  289.75,
  289.45,    289.45,  289.45,  289.45,
  289.15,    289.15,  289.15,  289.15,
  288.9,     288.9,   288.9,   288.9,
  288.35,    288.35,  288.35,  288.35,
  287.85,    287.85,  287.85,  287.85,
  287.7,     287.7,   287.7,   287.7,
  287.55,    287.55,  287.55,  287.55,
  287.35,    287.35,  287.35,  287.35,
  287.25,    287.25,  287.25,  287.25,
  287.55,    287.55,  287.55,  287.55,
  288.3,     288.3,   288.3,   288.3,
  289.1,     289.1,   289.1,   289.1,
  289.85,    289.85,  289.85,  289.85,
  290.5,     290.5,   290.5,   290.5,
  292.05,    292.05,  292.05,  292.05,
  294,       294,     294,     294,
  294.95,    294.95,  294.95,  294.95,
  295.35,    295.35,  295.35,  295.35,
  295.8,     295.8,   295.8,   295.8,
  295.95,    295.95,  295.95,  295.95,
  295.7,     295.7,   295.7,   295.7,
  295.9,     295.9,   295.9,   295.9,
  296.5,     296.5,   296.5,   296.5,
  297,       297,     297,     297,
  297.25,    297.25,  297.25,  297.25,
  297.55,    297.55,  297.55,  297.55,
  297.8,     297.8,   297.8,   297.8,
  298.15,    298.15,  298.15,  298.15,
  298.3,     298.3,   298.3,   298.3,
  298.25,    298.25,  298.25,  298.25,
  298.15,    298.15,  298.15,  298.15,
  297.5,     297.5,   297.5,   297.5,
  296.7,     296.7,   296.7,   296.7,
  296.2,     296.2,   296.2,   296.2,
  295.25,    295.25,  295.25,  295.25,
  292.6,     292.6,   292.6,   292.6,
  290.45,    290.45,  290.45,  290.45,
  290.1,     290.1,   290.1,   290.1,
  290,       290,     290,     290,
  289.85,    289.85,  289.85,  289.85,
  289.6,     289.6,   289.6,   289.6,
  289.45,    289.45,  289.45,  289.45,
  289.55,    289.55,  289.55,  289.55,
  289.75,    289.75,  289.75,  289.75,
  289.8,     289.8,   289.8,   289.8,
  289.55,    289.55,  289.55,  289.55,
  289.75,    289.75,  289.75,  289.75,
  289.55,    289.55,  289.55,  289.55,
  288.55,    288.55,  288.55,  288.55,
  288.2,     288.2,   288.2,   288.2,
  288.35,    288.35,  288.35,  288.35,
  288.1,     288.1,   288.1,   288.1,
  287.9,     287.9,   287.9,   287.9,
  288.1,     288.1,   288.1,   288.1,
  288.2,     288.2,   288.2,   288.2,
  288.25,    288.25,  288.25,  288.25,
  288.15,    288.15,  288.15,  288.15,
  288.25,    288.25,  288.25,  288.25,
  289,       289,     289,     289,
  289.85,    289.85,  289.85,  289.85,
  290.55,    290.55,  290.55,  290.55,
  291.35,    291.35,  291.35,  291.35,
  292.05,    292.05,  292.05,  292.05,
  292.8,     292.8,   292.8,   292.8,
  293.45,    293.45,  293.45,  293.45,
  293.4,     293.4,   293.4,   293.4,
  292.8,     292.8,   292.8,   292.8,
  292.5,     292.5,   292.5,   292.5,
  292.75,    292.75,  292.75,  292.75,
  293.15,    293.15,  293.15,  293.15,
  293.75,    293.75,  293.75,  293.75,
  294.35,    294.35,  294.35,  294.35,
  294.7,     294.7,   294.7,   294.7,
  294.95,    294.95,  294.95,  294.95,
  295.15,    295.15,  295.15,  295.15,
  295.15,    295.15,  295.15,  295.15,
  295.25,    295.25,  295.25,  295.25,
  295.5,     295.5,   295.5,   295.5,
  295.35,    295.35,  295.35,  295.35,
  295,       295,     295,     295,
  294.55,    294.55,  294.55,  294.55,
  294.1,     294.1,   294.1,   294.1,
  293.9,     293.9,   293.9,   293.9,
  293.55,    293.55,  293.55,  293.55,
  292.9,     292.9,   292.9,   292.9,
  292.05,    292.05,  292.05,  292.05,
  291.1,     291.1,   291.1,   291.1,
  290.25,    290.25,  290.25,  290.25,
  289.55,    289.55,  289.55,  289.55,
  289.15,    289.15,  289.15,  289.15,
  288.75,    288.75,  288.75,  288.75,
  288.15,    288.15,  288.15,  288.15,
  287.65,    287.65,  287.65,  287.65,
  287.55,    287.55,  287.55,  287.55,
  287.65,    287.65,  287.65,  287.65,
  287.6,     287.6,   287.6,   287.6,
  287.3,     287.3,   287.3,   287.3,
  286.85,    286.85,  286.85,  286.85,
  286.7,     286.7,   286.7,   286.7,
  286.6,     286.6,   286.6,   286.6,
  286.35,    286.35,  286.35,  286.35,
  286.15,    286.15,  286.15,  286.15,
  286.1,     286.1,   286.1,   286.1,
  286.05,    286.05,  286.05,  286.05,
  285.9,     285.9,   285.9,   285.9,
  286,       286,     286,     286,
  286.35,    286.35,  286.35,  286.35,
  286.8,     286.8,   286.8,   286.8,
  287.5,     287.5,   287.5,   287.5,
  288.35,    288.35,  288.35,  288.35,
  289.25,    289.25,  289.25,  289.25,
  290.25,    290.25,  290.25,  290.25,
  291.2,     291.2,   291.2,   291.2,
  291.8,     291.8,   291.8,   291.8,
  291.9,     291.9,   291.9,   291.9,
  291.95,    291.95,  291.95,  291.95,
  292.25,    292.25,  292.25,  292.25,
  292.1,     292.1,   292.1,   292.1,
  291.8,     291.8,   291.8,   291.8,
  291.95,    291.95,  291.95,  291.95,
  292.05,    292.05,  292.05,  292.05,
  292.15,    292.15,  292.15,  292.15,
  292.85,    292.85,  292.85,  292.85,
  293.75,    293.75,  293.75,  293.75,
  294.1,     294.1,   294.1,   294.1,
  293.3,     293.3,   293.3,   293.3,
  291.4,     291.4,   291.4,   291.4,
  290.2,     290.2,   290.2,   290.2,
  290.2,     290.2,   290.2,   290.2,
  290.7,     290.7,   290.7,   290.7,
  291.5,     291.5,   291.5,   291.5,
  291.8,     291.8,   291.8,   291.8,
  291.35,    291.35,  291.35,  291.35,
  290.9,     290.9,   290.9,   290.9,
  290.65,    290.65,  290.65,  290.65,
  290.65,    290.65,  290.65,  290.65,
  290.5,     290.5,   290.5,   290.5,
  289.6,     289.6,   289.6,   289.6,
  288.8,     288.8,   288.8,   288.8,
  288.45,    288.45,  288.45,  288.45,
  288,       288,     288,     288,
  287.5,     287.5,   287.5,   287.5,
  287.1,     287.1,   287.1,   287.1,
  287,       287,     287,     287,
  287.15,    287.15,  287.15,  287.15,
  287.3,     287.3,   287.3,   287.3,
  287.45,    287.45,  287.45,  287.45,
  287.65,    287.65,  287.65,  287.65,
  287.85,    287.85,  287.85,  287.85,
  287.95,    287.95,  287.95,  287.95,
  287.85,    287.85,  287.85,  287.85,
  287.7,     287.7,   287.7,   287.7,
  287.65,    287.65,  287.65,  287.65,
  287.8,     287.8,   287.8,   287.8,
  288.15,    288.15,  288.15,  288.15,
  288.6,     288.6,   288.6,   288.6,
  289.2,     289.2,   289.2,   289.2,
  289.8,     289.8,   289.8,   289.8,
  290.15,    290.15,  290.15,  290.15,
  290.15,    290.15,  290.15,  290.15,
  289.95,    289.95,  289.95,  289.95,
  289.9,     289.9,   289.9,   289.9,
  290.3,     290.3,   290.3,   290.3,
  291.35,    291.35,  291.35,  291.35,
  291.75,    291.75,  291.75,  291.75,
  291.5,     291.5,   291.5,   291.5,
  291.85,    291.85,  291.85,  291.85,
  292.35,    292.35,  292.35,  292.35,
  292.6,     292.6,   292.6,   292.6,
  292.6,     292.6,   292.6,   292.6,
  292.75,    292.75,  292.75,  292.75,
  293.2,     293.2,   293.2,   293.2,
  293.3,     293.3,   293.3,   293.3,
  293.1,     293.1,   293.1,   293.1,
  292.9,     292.9,   292.9,   292.9,
  292.6,     292.6,   292.6,   292.6,
  292.2,     292.2,   292.2,   292.2,
  291.85,    291.85,  291.85,  291.85,
  291.75,    291.75,  291.75,  291.75,
  291.4,     291.4,   291.4,   291.4,
  290.95,    290.95,  290.95,  290.95,
  290.7,     290.7,   290.7,   290.7,
  290.4,     290.4,   290.4,   290.4,
  290.15,    290.15,  290.15,  290.15,
  289.95,    289.95,  289.95,  289.95,
  289.8,     289.8,   289.8,   289.8,
  289.6,     289.6,   289.6,   289.6,
  289.4,     289.4,   289.4,   289.4,
  289.25,    289.25,  289.25,  289.25,
  289.15,    289.15,  289.15,  289.15,
  289.1,     289.1,   289.1,   289.1,
  289,       289,     289,     289,
  288.9,     288.9,   288.9,   288.9,
  288.8,     288.8,   288.8,   288.8,
  288.75,    288.75,  288.75,  288.75,
  288.7,     288.7,   288.7,   288.7,
  288.6,     288.6,   288.6,   288.6,
  288.5,     288.5,   288.5,   288.5,
  288.5,     288.5,   288.5,   288.5,
  288.5,     288.5,   288.5,   288.5,
  288.55,    288.55,  288.55,  288.55,
  288.8,     288.8,   288.8,   288.8,
  289.2,     289.2,   289.2,   289.2,
  289.65,    289.65,  289.65,  289.65,
  289.95,    289.95,  289.95,  289.95,
  290.3,     290.3,   290.3,   290.3,
  290.8,     290.8,   290.8,   290.8,
  291.4,     291.4,   291.4,   291.4,
  291.65,    291.65,  291.65,  291.65,
  291.5,     291.5,   291.5,   291.5,
  291.7,     291.7,   291.7,   291.7,
  291.75,    291.75,  291.75,  291.75,
  291.85,    291.85,  291.85,  291.85,
  292.35,    292.35,  292.35,  292.35,
  292.55,    292.55,  292.55,  292.55,
  292.45,    292.45,  292.45,  292.45,
  292.45,    292.45,  292.45,  292.45,
  292.6,     292.6,   292.6,   292.6,
  292.3,     292.3,   292.3,   292.3,
  291.75,    291.75,  291.75,  291.75,
  291.1,     291.1,   291.1,   291.1,
  290.5,     290.5,   290.5,   290.5,
  289.9,     289.9,   289.9,   289.9,
  289.05,    289.05,  289.05,  289.05,
  288.35,    288.35,  288.35,  288.35,
  288,       288,     288,     288,
  287.95,    287.95,  287.95,  287.95,
  288,       288,     288,     288,
  288.05,    288.05,  288.05,  288.05,
  288,       288,     288,     288,
  287.8,     287.8,   287.8,   287.8,
  287.5,     287.5,   287.5,   287.5,
  287.2,     287.2,   287.2,   287.2,
  286.75,    286.75,  286.75,  286.75,
  286.45,    286.45,  286.45,  286.45,
  286.45,    286.45,  286.45,  286.45,
  286.45,    286.45,  286.45,  286.45,
  286.4,     286.4,   286.4,   286.4,
  286.35,    286.35,  286.35,  286.35,
  286.35,    286.35,  286.35,  286.35,
  286.3,     286.3,   286.3,   286.3,
  286.25,    286.25,  286.25,  286.25,
  286.2,     286.2,   286.2,   286.2,
  286.1,     286.1,   286.1,   286.1,
  286,       286,     286,     286,
  285.95,    285.95,  285.95,  285.95,
  285.95,    285.95,  285.95,  285.95,
  285.9,     285.9,   285.9,   285.9,
  285.85,    285.85,  285.85,  285.85,
  286,       286,     286,     286,
  286.35,    286.35,  286.35,  286.35,
  286.85,    286.85,  286.85,  286.85,
  287.35,    287.35,  287.35,  287.35,
  287.65,    287.65,  287.65,  287.65,
  287.9,     287.9,   287.9,   287.9,
  288.2,     288.2,   288.2,   288.2,
  288.55,    288.55,  288.55,  288.55,
  289.1,     289.1,   289.1,   289.1,
  289.8,     289.8,   289.8,   289.8,
  290.45,    290.45,  290.45,  290.45,
  291.15,    291.15,  291.15,  291.15,
  291.8,     291.8,   291.8,   291.8,
  292,       292,     292,     292,
  291.45,    291.45,  291.45,  291.45,
  291,       291,     291,     291,
  291.1,     291.1,   291.1,   291.1,
  291.4,     291.4,   291.4,   291.4,
  291.85,    291.85,  291.85,  291.85,
  291.6,     291.6,   291.6,   291.6,
  291.25,    291.25,  291.25,  291.25,
  291.15,    291.15,  291.15,  291.15,
  290.8,     290.8,   290.8,   290.8,
  290.55,    290.55,  290.55,  290.55,
  290.5,     290.5,   290.5,   290.5,
  290.35,    290.35,  290.35,  290.35,
  289.95,    289.95,  289.95,  289.95,
  289.8,     289.8,   289.8,   289.8,
  289.9,     289.9,   289.9,   289.9,
  289.95,    289.95,  289.95,  289.95,
  289.9,     289.9,   289.9,   289.9,
  289.75,    289.75,  289.75,  289.75,
  289.6,     289.6,   289.6,   289.6,
  289.4,     289.4,   289.4,   289.4,
  289,       289,     289,     289,
  288.5,     288.5,   288.5,   288.5,
  288.15,    288.15,  288.15,  288.15,
  288,       288,     288,     288,
  287.9,     287.9,   287.9,   287.9,
  287.8,     287.8,   287.8,   287.8,
  287.75,    287.75,  287.75,  287.75,
  287.7,     287.7,   287.7,   287.7,
  287.55,    287.55,  287.55,  287.55,
  287.45,    287.45,  287.45,  287.45,
  287.4,     287.4,   287.4,   287.4,
  287.3,     287.3,   287.3,   287.3,
  287.2,     287.2,   287.2,   287.2,
  287.15,    287.15,  287.15,  287.15,
  287.25,    287.25,  287.25,  287.25,
  287.75,    287.75,  287.75,  287.75,
  288.5,     288.5,   288.5,   288.5,
  289.1,     289.1,   289.1,   289.1,
  289.6,     289.6,   289.6,   289.6,
  290.4,     290.4,   290.4,   290.4,
  291.4,     291.4,   291.4,   291.4,
  292.15,    292.15,  292.15,  292.15,
  292.7,     292.7,   292.7,   292.7,
  293.35,    293.35,  293.35,  293.35,
  293.95,    293.95,  293.95,  293.95,
  294.1,     294.1,   294.1,   294.1,
  294.2,     294.2,   294.2,   294.2,
  294.25,    294.25,  294.25,  294.25,
  292,       292,     292,     292,
  290.05,    290.05,  290.05,  290.05,
  291.1,     291.1,   291.1,   291.1,
  292.6,     292.6,   292.6,   292.6,
  293.5,     293.5,   293.5,   293.5,
  293.65,    293.65,  293.65,  293.65,
  293.9,     293.9,   293.9,   293.9,
  294.25,    294.25,  294.25,  294.25,
  294.35,    294.35,  294.35,  294.35,
  294.2,     294.2,   294.2,   294.2,
  293.95,    293.95,  293.95,  293.95,
  293.75,    293.75,  293.75,  293.75,
  293.25,    293.25,  293.25,  293.25,
  292.9,     292.9,   292.9,   292.9,
  292.45,    292.45,  292.45,  292.45,
  290.65,    290.65,  290.65,  290.65,
  288.8,     288.8,   288.8,   288.8,
  288.1,     288.1,   288.1,   288.1,
  287.75,    287.75,  287.75,  287.75,
  287.45,    287.45,  287.45,  287.45,
  287.2,     287.2,   287.2,   287.2,
  287.25,    287.25,  287.25,  287.25,
  287.2,     287.2,   287.2,   287.2,
  287.1,     287.1,   287.1,   287.1,
  287.1,     287.1,   287.1,   287.1,
  287.05,    287.05,  287.05,  287.05,
  286.95,    286.95,  286.95,  286.95,
  286.85,    286.85,  286.85,  286.85,
  286.75,    286.75,  286.75,  286.75,
  286.6,     286.6,   286.6,   286.6,
  286.45,    286.45,  286.45,  286.45,
  286.3,     286.3,   286.3,   286.3,
  286.2,     286.2,   286.2,   286.2,
  286.2,     286.2,   286.2,   286.2,
  286.45,    286.45,  286.45,  286.45,
  286.95,    286.95,  286.95,  286.95,
  287.6,     287.6,   287.6,   287.6,
  288.25,    288.25,  288.25,  288.25,
  289.15,    289.15,  289.15,  289.15,
  290.05,    290.05,  290.05,  290.05,
  290.85,    290.85,  290.85,  290.85,
  291.9,     291.9,   291.9,   291.9,
  292.75,    292.75,  292.75,  292.75,
  293.25,    293.25,  293.25,  293.25,
  293.5,     293.5,   293.5,   293.5,
  293.85,    293.85,  293.85,  293.85,
  294.15,    294.15,  294.15,  294.15,
  292.4,     292.4,   292.4,   292.4,
  290.8,     290.8,   290.8,   290.8,
  290.6,     290.6,   290.6,   290.6,
  290.35,    290.35,  290.35,  290.35,
  291.2,     291.2,   291.2,   291.2,
  292.4,     292.4,   292.4,   292.4,
  291.85,    291.85,  291.85,  291.85,
  291.15,    291.15,  291.15,  291.15,
  291.5,     291.5,   291.5,   291.5,
  291.25,    291.25,  291.25,  291.25,
  291.4,     291.4,   291.4,   291.4,
  292.2,     292.2,   292.2,   292.2,
  292.4,     292.4,   292.4,   292.4,
  292.35,    292.35,  292.35,  292.35,
  292.4,     292.4,   292.4,   292.4,
  292.1,     292.1,   292.1,   292.1,
  291.45,    291.45,  291.45,  291.45,
  290.6,     290.6,   290.6,   290.6,
  289.95,    289.95,  289.95,  289.95,
  289.5,     289.5,   289.5,   289.5,
  289.05,    289.05,  289.05,  289.05,
  288.7,     288.7,   288.7,   288.7,
  288.6,     288.6,   288.6,   288.6,
  288.65,    288.65,  288.65,  288.65,
  288.7,     288.7,   288.7,   288.7,
  288.75,    288.75,  288.75,  288.75,
  288.65,    288.65,  288.65,  288.65,
  288.55,    288.55,  288.55,  288.55,
  288.65,    288.65,  288.65,  288.65,
  288.95,    288.95,  288.95,  288.95,
  289.15,    289.15,  289.15,  289.15,
  289.1,     289.1,   289.1,   289.1,
  289.1,     289.1,   289.1,   289.1,
  289.25,    289.25,  289.25,  289.25,
  289.4,     289.4,   289.4,   289.4,
  289.75,    289.75,  289.75,  289.75,
  290.15,    290.15,  290.15,  290.15,
  290.4,     290.4,   290.4,   290.4,
  290.7,     290.7,   290.7,   290.7,
  291.3,     291.3,   291.3,   291.3,
  292.15,    292.15,  292.15,  292.15,
  292.8,     292.8,   292.8,   292.8,
  292.95,    292.95,  292.95,  292.95,
  293.4,     293.4,   293.4,   293.4,
  294.05,    294.05,  294.05,  294.05,
  294.1,     294.1,   294.1,   294.1,
  294.05,    294.05,  294.05,  294.05,
  294.1,     294.1,   294.1,   294.1,
  294.35,    294.35,  294.35,  294.35,
  294.6,     294.6,   294.6,   294.6,
  294.25,    294.25,  294.25,  294.25,
  293.45,    293.45,  293.45,  293.45,
  291.5,     291.5,   291.5,   291.5,
  289.95,    289.95,  289.95,  289.95,
  290.15,    290.15,  290.15,  290.15,
  290.2,     290.2,   290.2,   290.2,
  290.05,    290.05,  290.05,  290.05,
  290.1,     290.1,   290.1,   290.1,
  290.15,    290.15,  290.15,  290.15,
  290.15,    290.15,  290.15,  290.15,
  290.05,    290.05,  290.05,  290.05,
  289.9,     289.9,   289.9,   289.9,
  289.85,    289.85,  289.85,  289.85,
  289.85,    289.85,  289.85,  289.85,
  289.9,     289.9,   289.9,   289.9,
  290,       290,     290,     290,
  290.1,     290.1,   290.1,   290.1,
  290.2,     290.2,   290.2,   290.2,
  290.25,    290.25,  290.25,  290.25,
  290.25,    290.25,  290.25,  290.25,
  290.25,    290.25,  290.25,  290.25,
  290.25,    290.25,  290.25,  290.25,
  290.3,     290.3,   290.3,   290.3,
  290.35,    290.35,  290.35,  290.35,
  290.3,     290.3,   290.3,   290.3,
  290.25,    290.25,  290.25,  290.25,
  290.15,    290.15,  290.15,  290.15,
  289.9,     289.9,   289.9,   289.9,
  289.6,     289.6,   289.6,   289.6,
  289.35,    289.35,  289.35,  289.35,
  289.15,    289.15,  289.15,  289.15,
  288.95,    288.95,  288.95,  288.95,
  288.95,    288.95,  288.95,  288.95,
  289.05,    289.05,  289.05,  289.05,
  289.15,    289.15,  289.15,  289.15,
  289.3,     289.3,   289.3,   289.3,
  289.55,    289.55,  289.55,  289.55,
  289.85,    289.85,  289.85,  289.85,
  290.1,     290.1,   290.1,   290.1,
  290.5,     290.5,   290.5,   290.5,
  290.95,    290.95,  290.95,  290.95,
  291.2,     291.2,   291.2,   291.2,
  291.45,    291.45,  291.45,  291.45,
  292.05,    292.05,  292.05,  292.05,
  292.85,    292.85,  292.85,  292.85,
  293.5,     293.5,   293.5,   293.5,
  293.95,    293.95,  293.95,  293.95,
  294.2,     294.2,   294.2,   294.2,
  294.1,     294.1,   294.1,   294.1,
  293.65,    293.65,  293.65,  293.65,
  293.3,     293.3,   293.3,   293.3,
  293.55,    293.55,  293.55,  293.55,
  294.1,     294.1,   294.1,   294.1,
  294.1,     294.1,   294.1,   294.1,
  294,       294,     294,     294,
  294.4,     294.4,   294.4,   294.4,
  294.3,     294.3,   294.3,   294.3,
  293.85,    293.85,  293.85,  293.85,
  293.45,    293.45,  293.45,  293.45,
  293,       293,     293,     293,
  292.65,    292.65,  292.65,  292.65,
  292.1,     292.1,   292.1,   292.1,
  291.4,     291.4,   291.4,   291.4,
  290.95,    290.95,  290.95,  290.95,
  290.5,     290.5,   290.5,   290.5,
  289.85,    289.85,  289.85,  289.85,
  289.35,    289.35,  289.35,  289.35,
  288.95,    288.95,  288.95,  288.95,
  288.6,     288.6,   288.6,   288.6,
  288.45,    288.45,  288.45,  288.45,
  288.35,    288.35,  288.35,  288.35,
  288.1,     288.1,   288.1,   288.1,
  287.65,    287.65,  287.65,  287.65,
  287.05,    287.05,  287.05,  287.05,
  286.9,     286.9,   286.9,   286.9,
  287.2,     287.2,   287.2,   287.2,
  287.4,     287.4,   287.4,   287.4,
  287.55,    287.55,  287.55,  287.55,
  287.7,     287.7,   287.7,   287.7,
  287.75,    287.75,  287.75,  287.75,
  287.55,    287.55,  287.55,  287.55,
  287.35,    287.35,  287.35,  287.35,
  287.55,    287.55,  287.55,  287.55,
  288.05,    288.05,  288.05,  288.05,
  288.9,     288.9,   288.9,   288.9,
  289.95,    289.95,  289.95,  289.95,
  290.65,    290.65,  290.65,  290.65,
  291.05,    291.05,  291.05,  291.05,
  291.35,    291.35,  291.35,  291.35,
  291.75,    291.75,  291.75,  291.75,
  292.4,     292.4,   292.4,   292.4,
  292.95,    292.95,  292.95,  292.95,
  293.35,    293.35,  293.35,  293.35,
  293.9,     293.9,   293.9,   293.9,
  294.4,     294.4,   294.4,   294.4,
  294.55,    294.55,  294.55,  294.55,
  294.6,     294.6,   294.6,   294.6,
  295,       295,     295,     295,
  295.35,    295.35,  295.35,  295.35,
  295.55,    295.55,  295.55,  295.55,
  295.85,    295.85,  295.85,  295.85,
  295.95,    295.95,  295.95,  295.95,
  296.1,     296.1,   296.1,   296.1,
  296.15,    296.15,  296.15,  296.15,
  296,       296,     296,     296,
  295.9,     295.9,   295.9,   295.9,
  295.8,     295.8,   295.8,   295.8,
  295.55,    295.55,  295.55,  295.55,
  294.95,    294.95,  294.95,  294.95,
  294.2,     294.2,   294.2,   294.2,
  293.4,     293.4,   293.4,   293.4,
  292.65,    292.65,  292.65,  292.65,
  291.75,    291.75,  291.75,  291.75,
  290.8,     290.8,   290.8,   290.8,
  290.15,    290.15,  290.15,  290.15,
  289.55,    289.55,  289.55,  289.55,
  289.4,     289.4,   289.4,   289.4,
  289.45,    289.45,  289.45,  289.45,
  288.8,     288.8,   288.8,   288.8,
  288.25,    288.25,  288.25,  288.25,
  288.15,    288.15,  288.15,  288.15,
  288.25,    288.25,  288.25,  288.25,
  288.3,     288.3,   288.3,   288.3,
  287.95,    287.95,  287.95,  287.95,
  287.4,     287.4,   287.4,   287.4,
  286.8,     286.8,   286.8,   286.8,
  286.5,     286.5,   286.5,   286.5,
  286.5,     286.5,   286.5,   286.5,
  286.6,     286.6,   286.6,   286.6,
  286.85,    286.85,  286.85,  286.85,
  287.65,    287.65,  287.65,  287.65,
  289.1,     289.1,   289.1,   289.1,
  290.7,     290.7,   290.7,   290.7,
  291.8,     291.8,   291.8,   291.8,
  292.4,     292.4,   292.4,   292.4,
  292.85,    292.85,  292.85,  292.85,
  293.25,    293.25,  293.25,  293.25,
  293.7,     293.7,   293.7,   293.7,
  294.15,    294.15,  294.15,  294.15,
  294.5,     294.5,   294.5,   294.5,
  294.7,     294.7,   294.7,   294.7,
  294.75,    294.75,  294.75,  294.75,
  294.55,    294.55,  294.55,  294.55,
  293.3,     293.3,   293.3,   293.3,
  291.65,    291.65,  291.65,  291.65,
  290.8,     290.8,   290.8,   290.8,
  290.8,     290.8,   290.8,   290.8,
  291.1,     291.1,   291.1,   291.1,
  291.3,     291.3,   291.3,   291.3,
  291.8,     291.8,   291.8,   291.8,
  292.45,    292.45,  292.45,  292.45,
  293.2,     293.2,   293.2,   293.2,
  293.75,    293.75,  293.75,  293.75,
  293.75,    293.75,  293.75,  293.75,
  293.55,    293.55,  293.55,  293.55,
  293.3,     293.3,   293.3,   293.3,
  293,       293,     293,     293,
  292.7,     292.7,   292.7,   292.7,
  292.45,    292.45,  292.45,  292.45,
  292.25,    292.25,  292.25,  292.25,
  291.95,    291.95,  291.95,  291.95,
  291.45,    291.45,  291.45,  291.45,
  291,       291,     291,     291,
  290.3,     290.3,   290.3,   290.3,
  289.5,     289.5,   289.5,   289.5,
  289.25,    289.25,  289.25,  289.25,
  288.95,    288.95,  288.95,  288.95,
  288.75,    288.75,  288.75,  288.75,
  288.7,     288.7,   288.7,   288.7,
  288.55,    288.55,  288.55,  288.55,
  288.65,    288.65,  288.65,  288.65,
  288.75,    288.75,  288.75,  288.75,
  288.9,     288.9,   288.9,   288.9,
  289,       289,     289,     289,
  288.9,     288.9,   288.9,   288.9,
  288.7,     288.7,   288.7,   288.7,
  288.3,     288.3,   288.3,   288.3,
  287.95,    287.95,  287.95,  287.95,
  287.8,     287.8,   287.8,   287.8,
  287.65,    287.65,  287.65,  287.65,
  287.65,    287.65,  287.65,  287.65,
  287.95,    287.95,  287.95,  287.95,
  288.25,    288.25,  288.25,  288.25,
  288.2,     288.2,   288.2,   288.2,
  288.1,     288.1,   288.1,   288.1,
  288.45,    288.45,  288.45,  288.45,
  289.1,     289.1,   289.1,   289.1,
  290,       290,     290,     290,
  290.75,    290.75,  290.75,  290.75,
  290.6,     290.6,   290.6,   290.6,
  290.55,    290.55,  290.55,  290.55,
  290.75,    290.75,  290.75,  290.75,
  289.75,    289.75,  289.75,  289.75,
  289.6,     289.6,   289.6,   289.6,
  290.65,    290.65,  290.65,  290.65,
  291,       291,     291,     291,
  290.9,     290.9,   290.9,   290.9,
  290.5,     290.5,   290.5,   290.5,
  290,       290,     290,     290,
  289.55,    289.55,  289.55,  289.55,
  289.4,     289.4,   289.4,   289.4,
  289.7,     289.7,   289.7,   289.7,
  289.95,    289.95,  289.95,  289.95,
  289.9,     289.9,   289.9,   289.9,
  289.8,     289.8,   289.8,   289.8,
  289.55,    289.55,  289.55,  289.55,
  289.25,    289.25,  289.25,  289.25,
  288.9,     288.9,   288.9,   288.9,
  288.4,     288.4,   288.4,   288.4,
  287.95,    287.95,  287.95,  287.95,
  287.55,    287.55,  287.55,  287.55,
  287.3,     287.3,   287.3,   287.3,
  287.2,     287.2,   287.2,   287.2,
  287.25,    287.25,  287.25,  287.25,
  287.4,     287.4,   287.4,   287.4,
  287.65,    287.65,  287.65,  287.65,
  287.95,    287.95,  287.95,  287.95,
  288.1,     288.1,   288.1,   288.1,
  288.2,     288.2,   288.2,   288.2,
  288.3,     288.3,   288.3,   288.3,
  288.4,     288.4,   288.4,   288.4,
  288.45,    288.45,  288.45,  288.45,
  288.45,    288.45,  288.45,  288.45,
  288.4,     288.4,   288.4,   288.4,
  288.35,    288.35,  288.35,  288.35,
  288.5,     288.5,   288.5,   288.5,
  288.8,     288.8,   288.8,   288.8,
  289.1,     289.1,   289.1,   289.1,
  289.35,    289.35,  289.35,  289.35,
  289.8,     289.8,   289.8,   289.8,
  290.35,    290.35,  290.35,  290.35,
  290.7,     290.7,   290.7,   290.7,
  291.2,     291.2,   291.2,   291.2,
  291.85,    291.85,  291.85,  291.85,
  292.35,    292.35,  292.35,  292.35,
  292.75,    292.75,  292.75,  292.75,
  293.05,    293.05,  293.05,  293.05,
  293.4,     293.4,   293.4,   293.4,
  293.9,     293.9,   293.9,   293.9,
  294.4,     294.4,   294.4,   294.4,
  294.7,     294.7,   294.7,   294.7,
  294.55,    294.55,  294.55,  294.55,
  294.6,     294.6,   294.6,   294.6,
  294.85,    294.85,  294.85,  294.85,
  294.9,     294.9,   294.9,   294.9,
  294.95,    294.95,  294.95,  294.95,
  294.75,    294.75,  294.75,  294.75,
  294.5,     294.5,   294.5,   294.5,
  294.35,    294.35,  294.35,  294.35,
  294,       294,     294,     294,
  293.45,    293.45,  293.45,  293.45,
  293.1,     293.1,   293.1,   293.1,
  292.8,     292.8,   292.8,   292.8,
  292.3,     292.3,   292.3,   292.3,
  292,       292,     292,     292,
  291.7,     291.7,   291.7,   291.7,
  291.35,    291.35,  291.35,  291.35,
  290.8,     290.8,   290.8,   290.8,
  289.95,    289.95,  289.95,  289.95,
  289.6,     289.6,   289.6,   289.6,
  289.75,    289.75,  289.75,  289.75,
  290,       290,     290,     290,
  290.25,    290.25,  290.25,  290.25,
  290.5,     290.5,   290.5,   290.5,
  290.7,     290.7,   290.7,   290.7,
  290.95,    290.95,  290.95,  290.95,
  291.2,     291.2,   291.2,   291.2,
  291.15,    291.15,  291.15,  291.15,
  290.9,     290.9,   290.9,   290.9,
  290.75,    290.75,  290.75,  290.75,
  290.7,     290.7,   290.7,   290.7,
  290.7,     290.7,   290.7,   290.7,
  290.5,     290.5,   290.5,   290.5,
  290.15,    290.15,  290.15,  290.15,
  290.05,    290.05,  290.05,  290.05,
  290.05,    290.05,  290.05,  290.05,
  290.15,    290.15,  290.15,  290.15,
  290.5,     290.5,   290.5,   290.5,
  291,       291,     291,     291,
  291.4,     291.4,   291.4,   291.4,
  291.2,     291.2,   291.2,   291.2,
  290.5,     290.5,   290.5,   290.5,
  290.4,     290.4,   290.4,   290.4,
  290.6,     290.6,   290.6,   290.6,
  290.7,     290.7,   290.7,   290.7,
  290.95,    290.95,  290.95,  290.95,
  290.9,     290.9,   290.9,   290.9,
  290.75,    290.75,  290.75,  290.75,
  290.75,    290.75,  290.75,  290.75,
  290.45,    290.45,  290.45,  290.45,
  290.2,     290.2,   290.2,   290.2,
  290.55,    290.55,  290.55,  290.55,
  290.95,    290.95,  290.95,  290.95,
  290.8,     290.8,   290.8,   290.8,
  290.6,     290.6,   290.6,   290.6,
  290.7,     290.7,   290.7,   290.7,
  290.8,     290.8,   290.8,   290.8,
  290.85,    290.85,  290.85,  290.85,
  290.75,    290.75,  290.75,  290.75,
  290.5,     290.5,   290.5,   290.5,
  290.05,    290.05,  290.05,  290.05,
  289.35,    289.35,  289.35,  289.35,
  288.6,     288.6,   288.6,   288.6,
  288,       288,     288,     288,
  287.55,    287.55,  287.55,  287.55,
  287.1,     287.1,   287.1,   287.1,
  286.7,     286.7,   286.7,   286.7,
  286.45,    286.45,  286.45,  286.45,
  286.05,    286.05,  286.05,  286.05,
  285.7,     285.7,   285.7,   285.7,
  285.45,    285.45,  285.45,  285.45,
  285.35,    285.35,  285.35,  285.35,
  285.5,     285.5,   285.5,   285.5,
  285.3,     285.3,   285.3,   285.3,
  284.65,    284.65,  284.65,  284.65,
  284.05,    284.05,  284.05,  284.05,
  283.55,    283.55,  283.55,  283.55,
  283.2,     283.2,   283.2,   283.2,
  283.2,     283.2,   283.2,   283.2,
  283.35,    283.35,  283.35,  283.35,
  283.4,     283.4,   283.4,   283.4,
  283.45,    283.45,  283.45,  283.45,
  284,       284,     284,     284,
  285.25,    285.25,  285.25,  285.25,
  286.8,     286.8,   286.8,   286.8,
  288.65,    288.65,  288.65,  288.65,
  290.3,     290.3,   290.3,   290.3,
  291.3,     291.3,   291.3,   291.3,
  292.05,    292.05,  292.05,  292.05,
  292.65,    292.65,  292.65,  292.65,
  293.25,    293.25,  293.25,  293.25,
  293.9,     293.9,   293.9,   293.9,
  294.45,    294.45,  294.45,  294.45,
  294.75,    294.75,  294.75,  294.75,
  294.9,     294.9,   294.9,   294.9,
  295,       295,     295,     295,
  295.05,    295.05,  295.05,  295.05,
  295.2,     295.2,   295.2,   295.2,
  295,       295,     295,     295,
  294.6,     294.6,   294.6,   294.6,
  294.8,     294.8,   294.8,   294.8,
  294.85,    294.85,  294.85,  294.85,
  294.75,    294.75,  294.75,  294.75,
  294.95,    294.95,  294.95,  294.95,
  294.95,    294.95,  294.95,  294.95,
  294.55,    294.55,  294.55,  294.55,
  294,       294,     294,     294,
  293.4,     293.4,   293.4,   293.4,
  292.6,     292.6,   292.6,   292.6,
  291.75,    291.75,  291.75,  291.75,
  291.05,    291.05,  291.05,  291.05,
  290.5,     290.5,   290.5,   290.5,
  290.05,    290.05,  290.05,  290.05,
  289.5,     289.5,   289.5,   289.5,
  288.95,    288.95,  288.95,  288.95,
  288.6,     288.6,   288.6,   288.6,
  288.25,    288.25,  288.25,  288.25,
  287.8,     287.8,   287.8,   287.8,
  287.6,     287.6,   287.6,   287.6,
  287,       287,     287,     287,
  286.05,    286.05,  286.05,  286.05,
  285.95,    285.95,  285.95,  285.95,
  286.15,    286.15,  286.15,  286.15,
  286.1,     286.1,   286.1,   286.1,
  285.95,    285.95,  285.95,  285.95,
  285.5,     285.5,   285.5,   285.5,
  284.7,     284.7,   284.7,   284.7,
  284.2,     284.2,   284.2,   284.2,
  284.3,     284.3,   284.3,   284.3,
  284.75,    284.75,  284.75,  284.75,
  285.75,    285.75,  285.75,  285.75,
  287.1,     287.1,   287.1,   287.1,
  288.5,     288.5,   288.5,   288.5,
  289.9,     289.9,   289.9,   289.9,
  291.05,    291.05,  291.05,  291.05,
  291.95,    291.95,  291.95,  291.95,
  292.7,     292.7,   292.7,   292.7,
  293.35,    293.35,  293.35,  293.35,
  293.9,     293.9,   293.9,   293.9,
  294.05,    294.05,  294.05,  294.05,
  294.3,     294.3,   294.3,   294.3,
  294.9,     294.9,   294.9,   294.9,
  295.25,    295.25,  295.25,  295.25,
  295.55,    295.55,  295.55,  295.55,
  295.8,     295.8,   295.8,   295.8,
  296,       296,     296,     296,
  296.3,     296.3,   296.3,   296.3,
  296.55,    296.55,  296.55,  296.55,
  296.7,     296.7,   296.7,   296.7,
  296.7,     296.7,   296.7,   296.7,
  296.75,    296.75,  296.75,  296.75,
  296.75,    296.75,  296.75,  296.75,
  296.65,    296.65,  296.65,  296.65,
  296.5,     296.5,   296.5,   296.5,
  296.35,    296.35,  296.35,  296.35,
  296.15,    296.15,  296.15,  296.15,
  295.7,     295.7,   295.7,   295.7,
  295.15,    295.15,  295.15,  295.15,
  294.35,    294.35,  294.35,  294.35,
  293.1,     293.1,   293.1,   293.1,
  292.05,    292.05,  292.05,  292.05,
  291.4,     291.4,   291.4,   291.4,
  290.8,     290.8,   290.8,   290.8,
  290.4,     290.4,   290.4,   290.4,
  290.2,     290.2,   290.2,   290.2,
  289.9,     289.9,   289.9,   289.9,
  289.35,    289.35,  289.35,  289.35,
  288.9,     288.9,   288.9,   288.9,
  288.55,    288.55,  288.55,  288.55,
  288.3,     288.3,   288.3,   288.3,
  288.15,    288.15,  288.15,  288.15,
  288.15,    288.15,  288.15,  288.15,
  288.25,    288.25,  288.25,  288.25,
  288.15,    288.15,  288.15,  288.15,
  287.95,    287.95,  287.95,  287.95,
  287.9,     287.9,   287.9,   287.9,
  288.15,    288.15,  288.15,  288.15,
  288.75,    288.75,  288.75,  288.75,
  289.5,     289.5,   289.5,   289.5,
  290.25,    290.25,  290.25,  290.25,
  291.1,     291.1,   291.1,   291.1,
  291.9,     291.9,   291.9,   291.9,
  292.65,    292.65,  292.65,  292.65,
  293.15,    293.15,  293.15,  293.15,
  293.55,    293.55,  293.55,  293.55,
  294.3,     294.3,   294.3,   294.3,
  295.3,     295.3,   295.3,   295.3,
  296.05,    296.05,  296.05,  296.05,
  296.35,    296.35,  296.35,  296.35,
  296.55,    296.55,  296.55,  296.55,
  296.65,    296.65,  296.65,  296.65,
  296.65,    296.65,  296.65,  296.65,
  296.4,     296.4,   296.4,   296.4,
  295.95,    295.95,  295.95,  295.95,
  295.35,    295.35,  295.35,  295.35,
  294.65,    294.65,  294.65,  294.65,
  294.15,    294.15,  294.15,  294.15,
  294.1,     294.1,   294.1,   294.1,
  294.25,    294.25,  294.25,  294.25,
  294.6,     294.6,   294.6,   294.6,
  294.95,    294.95,  294.95,  294.95,
  294.45,    294.45,  294.45,  294.45,
  293.65,    293.65,  293.65,  293.65,
  293.35,    293.35,  293.35,  293.35,
  292.8,     292.8,   292.8,   292.8,
  291.7,     291.7,   291.7,   291.7,
  290.65,    290.65,  290.65,  290.65,
  289.7,     289.7,   289.7,   289.7,
  289.1,     289.1,   289.1,   289.1,
  288.75,    288.75,  288.75,  288.75,
  288.4,     288.4,   288.4,   288.4,
  287.9,     287.9,   287.9,   287.9,
  287.3,     287.3,   287.3,   287.3,
  286.9,     286.9,   286.9,   286.9,
  286.75,    286.75,  286.75,  286.75,
  286.8,     286.8,   286.8,   286.8,
  286.9,     286.9,   286.9,   286.9,
  287,       287,     287,     287,
  287.05,    287.05,  287.05,  287.05,
  287.25,    287.25,  287.25,  287.25,
  287.5,     287.5,   287.5,   287.5,
  287.65,    287.65,  287.65,  287.65,
  287.75,    287.75,  287.75,  287.75,
  287.8,     287.8,   287.8,   287.8,
  287.85,    287.85,  287.85,  287.85,
  287.95,    287.95,  287.95,  287.95,
  288.3,     288.3,   288.3,   288.3,
  288.7,     288.7,   288.7,   288.7,
  289.1,     289.1,   289.1,   289.1,
  289.8,     289.8,   289.8,   289.8,
  290.25,    290.25,  290.25,  290.25,
  289.85,    289.85,  289.85,  289.85,
  288.7,     288.7,   288.7,   288.7,
  288.6,     288.6,   288.6,   288.6,
  289.75,    289.75,  289.75,  289.75,
  290.2,     290.2,   290.2,   290.2,
  290.25,    290.25,  290.25,  290.25,
  290.55,    290.55,  290.55,  290.55,
  290.9,     290.9,   290.9,   290.9,
  291.05,    291.05,  291.05,  291.05,
  291,       291,     291,     291,
  290.75,    290.75,  290.75,  290.75,
  289.35,    289.35,  289.35,  289.35,
  287.8,     287.8,   287.8,   287.8,
  287.65,    287.65,  287.65,  287.65,
  288.05,    288.05,  288.05,  288.05,
  288.5,     288.5,   288.5,   288.5,
  288.85,    288.85,  288.85,  288.85,
  289.1,     289.1,   289.1,   289.1,
  289.15,    289.15,  289.15,  289.15,
  289.05,    289.05,  289.05,  289.05,
  288.85,    288.85,  288.85,  288.85,
  288.5,     288.5,   288.5,   288.5,
  288.25,    288.25,  288.25,  288.25,
  288,       288,     288,     288,
  287.7,     287.7,   287.7,   287.7,
  287.2,     287.2,   287.2,   287.2,
  286.7,     286.7,   286.7,   286.7,
  286.55,    286.55,  286.55,  286.55,
  286.55,    286.55,  286.55,  286.55,
  286.55,    286.55,  286.55,  286.55,
  286.55,    286.55,  286.55,  286.55,
  286.55,    286.55,  286.55,  286.55,
  286.6,     286.6,   286.6,   286.6,
  286.65,    286.65,  286.65,  286.65,
  286.65,    286.65,  286.65,  286.65,
  286.65,    286.65,  286.65,  286.65,
  286.7,     286.7,   286.7,   286.7,
  286.75,    286.75,  286.75,  286.75,
  286.75,    286.75,  286.75,  286.75,
  286.75,    286.75,  286.75,  286.75,
  286.75,    286.75,  286.75,  286.75,
  286.75,    286.75,  286.75,  286.75,
  286.8,     286.8,   286.8,   286.8,
  286.9,     286.9,   286.9,   286.9,
  287.05,    287.05,  287.05,  287.05,
  287.25,    287.25,  287.25,  287.25,
  287.5,     287.5,   287.5,   287.5,
  287.85,    287.85,  287.85,  287.85,
  288.1,     288.1,   288.1,   288.1,
  288.15,    288.15,  288.15,  288.15,
  288.25,    288.25,  288.25,  288.25,
  288.8,     288.8,   288.8,   288.8,
  289.65,    289.65,  289.65,  289.65,
  290.3,     290.3,   290.3,   290.3,
  290.7,     290.7,   290.7,   290.7,
  291.2,     291.2,   291.2,   291.2,
  291.9,     291.9,   291.9,   291.9,
  292.2,     292.2,   292.2,   292.2,
  292.3,     292.3,   292.3,   292.3,
  292.5,     292.5,   292.5,   292.5,
  292.55,    292.55,  292.55,  292.55,
  292.6,     292.6,   292.6,   292.6,
  292.6,     292.6,   292.6,   292.6,
  292.35,    292.35,  292.35,  292.35,
  292,       292,     292,     292,
  291.8,     291.8,   291.8,   291.8,
  291.6,     291.6,   291.6,   291.6,
  291.35,    291.35,  291.35,  291.35,
  291.1,     291.1,   291.1,   291.1,
  290.8,     290.8,   290.8,   290.8,
  290.45,    290.45,  290.45,  290.45,
  289.9,     289.9,   289.9,   289.9,
  289.4,     289.4,   289.4,   289.4,
  289.2,     289.2,   289.2,   289.2,
  289.1,     289.1,   289.1,   289.1,
  289,       289,     289,     289,
  288.9,     288.9,   288.9,   288.9,
  288.85,    288.85,  288.85,  288.85,
  288.85,    288.85,  288.85,  288.85,
  288.9,     288.9,   288.9,   288.9,
  288.95,    288.95,  288.95,  288.95,
  289,       289,     289,     289,
  289.1,     289.1,   289.1,   289.1,
  289.2,     289.2,   289.2,   289.2,
  289.3,     289.3,   289.3,   289.3,
  289.4,     289.4,   289.4,   289.4,
  289.5,     289.5,   289.5,   289.5,
  289.55,    289.55,  289.55,  289.55,
  289.6,     289.6,   289.6,   289.6,
  289.75,    289.75,  289.75,  289.75,
  289.9,     289.9,   289.9,   289.9,
  290.05,    290.05,  290.05,  290.05,
  290.3,     290.3,   290.3,   290.3,
  290.5,     290.5,   290.5,   290.5,
  290.55,    290.55,  290.55,  290.55,
  290.6,     290.6,   290.6,   290.6,
  290.8,     290.8,   290.8,   290.8,
  291.45,    291.45,  291.45,  291.45,
  292.15,    292.15,  292.15,  292.15,
  292.75,    292.75,  292.75,  292.75,
  293.05,    293.05,  293.05,  293.05,
  293.25,    293.25,  293.25,  293.25,
  293.75,    293.75,  293.75,  293.75,
  294.1,     294.1,   294.1,   294.1,
  294.35,    294.35,  294.35,  294.35,
  294.5,     294.5,   294.5,   294.5,
  294.55,    294.55,  294.55,  294.55,
  294.65,    294.65,  294.65,  294.65,
  294.6,     294.6,   294.6,   294.6,
  294.35,    294.35,  294.35,  294.35,
  294.2,     294.2,   294.2,   294.2,
  294.15,    294.15,  294.15,  294.15,
  293.95,    293.95,  293.95,  293.95,
  293.7,     293.7,   293.7,   293.7,
  293.7,     293.7,   293.7,   293.7,
  293.45,    293.45,  293.45,  293.45,
  292.75,    292.75,  292.75,  292.75,
  292.2,     292.2,   292.2,   292.2,
  292.05,    292.05,  292.05,  292.05,
  291.9,     291.9,   291.9,   291.9,
  291.45,    291.45,  291.45,  291.45,
  290.6,     290.6,   290.6,   290.6,
  289.5,     289.5,   289.5,   289.5,
  288.85,    288.85,  288.85,  288.85,
  288.35,    288.35,  288.35,  288.35,
  287.7,     287.7,   287.7,   287.7,
  287.3,     287.3,   287.3,   287.3,
  287.25,    287.25,  287.25,  287.25,
  287.55,    287.55,  287.55,  287.55,
  287.65,    287.65,  287.65,  287.65,
  287.4,     287.4,   287.4,   287.4,
  287,       287,     287,     287,
  286.75,    286.75,  286.75,  286.75,
  286.75,    286.75,  286.75,  286.75,
  286.9,     286.9,   286.9,   286.9,
  287.05,    287.05,  287.05,  287.05,
  287,       287,     287,     287,
  287,       287,     287,     287,
  287.1,     287.1,   287.1,   287.1,
  287.45,    287.45,  287.45,  287.45,
  288,       288,     288,     288,
  288.5,     288.5,   288.5,   288.5,
  289.05,    289.05,  289.05,  289.05,
  289.75,    289.75,  289.75,  289.75,
  290.4,     290.4,   290.4,   290.4,
  290.8,     290.8,   290.8,   290.8,
  291.3,     291.3,   291.3,   291.3,
  291.75,    291.75,  291.75,  291.75,
  292.05,    292.05,  292.05,  292.05,
  292.4,     292.4,   292.4,   292.4,
  292.65,    292.65,  292.65,  292.65,
  292.85,    292.85,  292.85,  292.85,
  293.35,    293.35,  293.35,  293.35,
  293.7,     293.7,   293.7,   293.7,
  293.5,     293.5,   293.5,   293.5,
  293.55,    293.55,  293.55,  293.55,
  293.6,     293.6,   293.6,   293.6,
  293.4,     293.4,   293.4,   293.4,
  293.3,     293.3,   293.3,   293.3,
  293.2,     293.2,   293.2,   293.2,
  293.15,    293.15,  293.15,  293.15,
  293.05,    293.05,  293.05,  293.05,
  292.8,     292.8,   292.8,   292.8,
  292.5,     292.5,   292.5,   292.5,
  292.2,     292.2,   292.2,   292.2,
  291.95,    291.95,  291.95,  291.95,
  291.75,    291.75,  291.75,  291.75,
  291.55,    291.55,  291.55,  291.55,
  291.3,     291.3,   291.3,   291.3,
  290.95,    290.95,  290.95,  290.95,
  290.65,    290.65,  290.65,  290.65,
  290.55,    290.55,  290.55,  290.55,
  290.45,    290.45,  290.45,  290.45,
  290.25,    290.25,  290.25,  290.25,
  289.95,    289.95,  289.95,  289.95,
  289.6,     289.6,   289.6,   289.6,
  289.3,     289.3,   289.3,   289.3,
  289.1,     289.1,   289.1,   289.1,
  288.9,     288.9,   288.9,   288.9,
  288.55,    288.55,  288.55,  288.55,
  288.2,     288.2,   288.2,   288.2,
  287.9,     287.9,   287.9,   287.9,
  287.75,    287.75,  287.75,  287.75,
  287.9,     287.9,   287.9,   287.9,
  288,       288,     288,     288,
  287.95,    287.95,  287.95,  287.95,
  288.1,     288.1,   288.1,   288.1,
  288.55,    288.55,  288.55,  288.55,
  289.1,     289.1,   289.1,   289.1,
  289.45,    289.45,  289.45,  289.45,
  289.85,    289.85,  289.85,  289.85,
  290.4,     290.4,   290.4,   290.4,
  291.1,     291.1,   291.1,   291.1,
  291.8,     291.8,   291.8,   291.8,
  292.3,     292.3,   292.3,   292.3,
  292.6,     292.6,   292.6,   292.6,
  292.9,     292.9,   292.9,   292.9,
  293.4,     293.4,   293.4,   293.4,
  293.8,     293.8,   293.8,   293.8,
  294.25,    294.25,  294.25,  294.25,
  294.75,    294.75,  294.75,  294.75,
  295.15,    295.15,  295.15,  295.15,
  295.15,    295.15,  295.15,  295.15,
  294.85,    294.85,  294.85,  294.85,
  294.7,     294.7,   294.7,   294.7,
  294.7,     294.7,   294.7,   294.7,
  294.8,     294.8,   294.8,   294.8,
  294.75,    294.75,  294.75,  294.75,
  294.75,    294.75,  294.75,  294.75,
  294.75,    294.75,  294.75,  294.75,
  294.4,     294.4,   294.4,   294.4,
  293.95,    293.95,  293.95,  293.95,
  293.45,    293.45,  293.45,  293.45,
  292.8,     292.8,   292.8,   292.8,
  291.95,    291.95,  291.95,  291.95,
  291.05,    291.05,  291.05,  291.05,
  290.25,    290.25,  290.25,  290.25,
  289.45,    289.45,  289.45,  289.45,
  288.8,     288.8,   288.8,   288.8,
  288.35,    288.35,  288.35,  288.35,
  288.05,    288.05,  288.05,  288.05,
  287.85,    287.85,  287.85,  287.85,
  287.6,     287.6,   287.6,   287.6,
  287.3,     287.3,   287.3,   287.3,
  287,       287,     287,     287,
  286.65,    286.65,  286.65,  286.65,
  286.2,     286.2,   286.2,   286.2,
  285.65,    285.65,  285.65,  285.65,
  285.25,    285.25,  285.25,  285.25,
  285.1,     285.1,   285.1,   285.1,
  284.75,    284.75,  284.75,  284.75,
  284.1,     284.1,   284.1,   284.1,
  283.55,    283.55,  283.55,  283.55,
  283.45,    283.45,  283.45,  283.45,
  283.75,    283.75,  283.75,  283.75,
  284.15,    284.15,  284.15,  284.15,
  285,       285,     285,     285,
  286.6,     286.6,   286.6,   286.6,
  288,       288,     288,     288,
  288.95,    288.95,  288.95,  288.95,
  289.65,    289.65,  289.65,  289.65,
  290.05,    290.05,  290.05,  290.05,
  290.65,    290.65,  290.65,  290.65,
  291.2,     291.2,   291.2,   291.2,
  291.9,     291.9,   291.9,   291.9,
  292.75,    292.75,  292.75,  292.75,
  293.4,     293.4,   293.4,   293.4,
  294.05,    294.05,  294.05,  294.05,
  294.55,    294.55,  294.55,  294.55,
  295.05,    295.05,  295.05,  295.05,
  295.6,     295.6,   295.6,   295.6,
  296.2,     296.2,   296.2,   296.2,
  296.6,     296.6,   296.6,   296.6,
  296.65,    296.65,  296.65,  296.65,
  296.6,     296.6,   296.6,   296.6,
  297.05,    297.05,  297.05,  297.05,
  297.45,    297.45,  297.45,  297.45,
  297.3,     297.3,   297.3,   297.3,
  297.25,    297.25,  297.25,  297.25,
  296.85,    296.85,  296.85,  296.85,
  296.35,    296.35,  296.35,  296.35,
  295.75,    295.75,  295.75,  295.75,
  294.7,     294.7,   294.7,   294.7,
  293.65,    293.65,  293.65,  293.65,
  292.9,     292.9,   292.9,   292.9,
  292.5,     292.5,   292.5,   292.5,
  292.15,    292.15,  292.15,  292.15,
  291.85,    291.85,  291.85,  291.85,
  291.55,    291.55,  291.55,  291.55,
  291.2,     291.2,   291.2,   291.2,
  290.9,     290.9,   290.9,   290.9,
  290.7,     290.7,   290.7,   290.7,
  290.55,    290.55,  290.55,  290.55,
  290.4,     290.4,   290.4,   290.4,
  290.35,    290.35,  290.35,  290.35,
  290.3,     290.3,   290.3,   290.3,
  290.15,    290.15,  290.15,  290.15,
  289.95,    289.95,  289.95,  289.95,
  289.75,    289.75,  289.75,  289.75,
  289.45,    289.45,  289.45,  289.45,
  289.15,    289.15,  289.15,  289.15,
  288.95,    288.95,  288.95,  288.95,
  289.05,    289.05,  289.05,  289.05,
  289.6,     289.6,   289.6,   289.6,
  290.35,    290.35,  290.35,  290.35,
  291.25,    291.25,  291.25,  291.25,
  292.2,     292.2,   292.2,   292.2,
  293.1,     293.1,   293.1,   293.1,
  294.05,    294.05,  294.05,  294.05,
  295.15,    295.15,  295.15,  295.15,
  296.05,    296.05,  296.05,  296.05,
  296.6,     296.6,   296.6,   296.6,
  297.1,     297.1,   297.1,   297.1,
  297.55,    297.55,  297.55,  297.55,
  297.9,     297.9,   297.9,   297.9,
  298.25,    298.25,  298.25,  298.25,
  298.6,     298.6,   298.6,   298.6,
  298.75,    298.75,  298.75,  298.75,
  298.85,    298.85,  298.85,  298.85,
  299.05,    299.05,  299.05,  299.05,
  299.2,     299.2,   299.2,   299.2,
  299.15,    299.15,  299.15,  299.15,
  299.05,    299.05,  299.05,  299.05,
  299.1,     299.1,   299.1,   299.1,
  299.1,     299.1,   299.1,   299.1,
  298.95,    298.95,  298.95,  298.95,
  298.75,    298.75,  298.75,  298.75,
  298.45,    298.45,  298.45,  298.45,
  298,       298,     298,     298,
  297.4,     297.4,   297.4,   297.4,
  296.55,    296.55,  296.55,  296.55,
  295.55,    295.55,  295.55,  295.55,
  294.8,     294.8,   294.8,   294.8,
  294.35,    294.35,  294.35,  294.35,
  294.05,    294.05,  294.05,  294.05,
  293.95,    293.95,  293.95,  293.95,
  293.8,     293.8,   293.8,   293.8,
  293.45,    293.45,  293.45,  293.45,
  293,       293,     293,     293,
  292.55,    292.55,  292.55,  292.55,
  292.1,     292.1,   292.1,   292.1,
  291.65,    291.65,  291.65,  291.65,
  291.25,    291.25,  291.25,  291.25,
  291,       291,     291,     291,
  290.75,    290.75,  290.75,  290.75,
  290.4,     290.4,   290.4,   290.4,
  290.05,    290.05,  290.05,  290.05,
  289.7,     289.7,   289.7,   289.7,
  289.5,     289.5,   289.5,   289.5,
  289.5,     289.5,   289.5,   289.5,
  289.85,    289.85,  289.85,  289.85,
  290.6,     290.6,   290.6,   290.6,
  291.35,    291.35,  291.35,  291.35,
  291.9,     291.9,   291.9,   291.9,
  292.6,     292.6,   292.6,   292.6,
  293.6,     293.6,   293.6,   293.6,
  294.65,    294.65,  294.65,  294.65,
  295.4,     295.4,   295.4,   295.4,
  295.85,    295.85,  295.85,  295.85,
  296.4,     296.4,   296.4,   296.4,
  297.1,     297.1,   297.1,   297.1,
  297.65,    297.65,  297.65,  297.65,
  298.1,     298.1,   298.1,   298.1,
  298.5,     298.5,   298.5,   298.5,
  298.7,     298.7,   298.7,   298.7,
  298.75,    298.75,  298.75,  298.75,
  298.9,     298.9,   298.9,   298.9,
  299.15,    299.15,  299.15,  299.15,
  299.4,     299.4,   299.4,   299.4,
  299.5,     299.5,   299.5,   299.5,
  299.6,     299.6,   299.6,   299.6,
  299.6,     299.6,   299.6,   299.6,
  299.5,     299.5,   299.5,   299.5,
  299.35,    299.35,  299.35,  299.35,
  299.15,    299.15,  299.15,  299.15,
  299,       299,     299,     299,
  298.5,     298.5,   298.5,   298.5,
  297.8,     297.8,   297.8,   297.8,
  296.9,     296.9,   296.9,   296.9,
  295.9,     295.9,   295.9,   295.9,
  295.3,     295.3,   295.3,   295.3,
  294.9,     294.9,   294.9,   294.9,
  294.55,    294.55,  294.55,  294.55,
  294.3,     294.3,   294.3,   294.3,
  294,       294,     294,     294,
  293.75,    293.75,  293.75,  293.75,
  293.35,    293.35,  293.35,  293.35,
  292.75,    292.75,  292.75,  292.75,
  292.25,    292.25,  292.25,  292.25,
  291.9,     291.9,   291.9,   291.9,
  291.75,    291.75,  291.75,  291.75,
  291.7,     291.7,   291.7,   291.7,
  291.55,    291.55,  291.55,  291.55,
  291.3,     291.3,   291.3,   291.3,
  291.05,    291.05,  291.05,  291.05,
  290.9,     290.9,   290.9,   290.9,
  290.6,     290.6,   290.6,   290.6,
  290.25,    290.25,  290.25,  290.25,
  290.2,     290.2,   290.2,   290.2,
  290.6,     290.6,   290.6,   290.6,
  291.35,    291.35,  291.35,  291.35,
  292.2,     292.2,   292.2,   292.2,
  293.25,    293.25,  293.25,  293.25,
  294.5,     294.5,   294.5,   294.5,
  295.85,    295.85,  295.85,  295.85,
  296.85,    296.85,  296.85,  296.85,
  297.7,     297.7,   297.7,   297.7,
  298.45,    298.45,  298.45,  298.45,
  298.9,     298.9,   298.9,   298.9,
  299.25,    299.25,  299.25,  299.25,
  299.45,    299.45,  299.45,  299.45,
  299.75,    299.75,  299.75,  299.75,
  300.1,     300.1,   300.1,   300.1,
  300.2,     300.2,   300.2,   300.2,
  300.2,     300.2,   300.2,   300.2,
  300.4,     300.4,   300.4,   300.4,
  300.6,     300.6,   300.6,   300.6,
  300.5,     300.5,   300.5,   300.5,
  300.45,    300.45,  300.45,  300.45,
  300.65,    300.65,  300.65,  300.65,
  300.35,    300.35,  300.35,  300.35,
  300.05,    300.05,  300.05,  300.05,
  300.15,    300.15,  300.15,  300.15,
  299.95,    299.95,  299.95,  299.95,
  299.45,    299.45,  299.45,  299.45,
  298.75,    298.75,  298.75,  298.75,
  298,       298,     298,     298,
  297.05,    297.05,  297.05,  297.05,
  295.95,    295.95,  295.95,  295.95,
  295.3,     295.3,   295.3,   295.3,
  294.8,     294.8,   294.8,   294.8,
  294.1,     294.1,   294.1,   294.1,
  293.75,    293.75,  293.75,  293.75,
  293.5,     293.5,   293.5,   293.5,
  293.25,    293.25,  293.25,  293.25,
  293.2,     293.2,   293.2,   293.2,
  293.1,     293.1,   293.1,   293.1,
  292.95,    292.95,  292.95,  292.95,
  292.5,     292.5,   292.5,   292.5,
  292.1,     292.1,   292.1,   292.1,
  291.9,     291.9,   291.9,   291.9,
  291.45,    291.45,  291.45,  291.45,
  291,       291,     291,     291,
  290.7,     290.7,   290.7,   290.7,
  290.35,    290.35,  290.35,  290.35,
  290.2,     290.2,   290.2,   290.2,
  290.4,     290.4,   290.4,   290.4,
  291.1,     291.1,   291.1,   291.1,
  292.4,     292.4,   292.4,   292.4,
  293.9,     293.9,   293.9,   293.9,
  295.35,    295.35,  295.35,  295.35,
  296.75,    296.75,  296.75,  296.75,
  297.8,     297.8,   297.8,   297.8,
  298.75,    298.75,  298.75,  298.75,
  299.65,    299.65,  299.65,  299.65,
  300.05,    300.05,  300.05,  300.05,
  300.4,     300.4,   300.4,   300.4,
  300.5,     300.5,   300.5,   300.5,
  300.25,    300.25,  300.25,  300.25,
  300.25,    300.25,  300.25,  300.25,
  300.4,     300.4,   300.4,   300.4,
  300.5,     300.5,   300.5,   300.5,
  300.85,    300.85,  300.85,  300.85,
  301.5,     301.5,   301.5,   301.5,
  301.75,    301.75,  301.75,  301.75,
  301.55,    301.55,  301.55,  301.55,
  301.4,     301.4,   301.4,   301.4,
  301.2,     301.2,   301.2,   301.2,
  300.95,    300.95,  300.95,  300.95,
  300.7,     300.7,   300.7,   300.7,
  300.45,    300.45,  300.45,  300.45,
  300.05,    300.05,  300.05,  300.05,
  299.55,    299.55,  299.55,  299.55,
  298.9,     298.9,   298.9,   298.9,
  297.8,     297.8,   297.8,   297.8,
  296.85,    296.85,  296.85,  296.85,
  295.9,     295.9,   295.9,   295.9,
  295.25,    295.25,  295.25,  295.25,
  295.2,     295.2,   295.2,   295.2,
  294.7,     294.7,   294.7,   294.7,
  293.95,    293.95,  293.95,  293.95,
  293.45,    293.45,  293.45,  293.45,
  293.1,     293.1,   293.1,   293.1,
  292.95,    292.95,  292.95,  292.95,
  292.75,    292.75,  292.75,  292.75,
  292.45,    292.45,  292.45,  292.45,
  292.4,     292.4,   292.4,   292.4,
  292.35,    292.35,  292.35,  292.35,
  292.7,     292.7,   292.7,   292.7,
  292.8,     292.8,   292.8,   292.8,
  292.4,     292.4,   292.4,   292.4,
  292.2,     292.2,   292.2,   292.2,
  291.9,     291.9,   291.9,   291.9,
  292.05,    292.05,  292.05,  292.05,
  292.15,    292.15,  292.15,  292.15,
  291.8,     291.8,   291.8,   291.8,
  292.15,    292.15,  292.15,  292.15,
  293.5,     293.5,   293.5,   293.5,
  295.05,    295.05,  295.05,  295.05,
  296.35,    296.35,  296.35,  296.35,
  297.55,    297.55,  297.55,  297.55,
  298.8,     298.8,   298.8,   298.8,
  300.1,     300.1,   300.1,   300.1,
  301.2,     301.2,   301.2,   301.2,
  302,       302,     302,     302,
  302.4,     302.4,   302.4,   302.4,
  302.55,    302.55,  302.55,  302.55,
  302.7,     302.7,   302.7,   302.7,
  302.7,     302.7,   302.7,   302.7,
  302.65,    302.65,  302.65,  302.65,
  302.8,     302.8,   302.8,   302.8,
  302.95,    302.95,  302.95,  302.95,
  302.85,    302.85,  302.85,  302.85,
  302.75,    302.75,  302.75,  302.75,
  302.85,    302.85,  302.85,  302.85,
  302.9,     302.9,   302.9,   302.9,
  302.85,    302.85,  302.85,  302.85,
  302.75,    302.75,  302.75,  302.75,
  302.55,    302.55,  302.55,  302.55,
  302.25,    302.25,  302.25,  302.25,
  301.7,     301.7,   301.7,   301.7,
  300.85,    300.85,  300.85,  300.85,
  299.85,    299.85,  299.85,  299.85,
  298.95,    298.95,  298.95,  298.95,
  298.25,    298.25,  298.25,  298.25,
  297.75,    297.75,  297.75,  297.75,
  297.4,     297.4,   297.4,   297.4,
  297.2,     297.2,   297.2,   297.2,
  296.9,     296.9,   296.9,   296.9,
  296.3,     296.3,   296.3,   296.3,
  295.9,     295.9,   295.9,   295.9,
  295.8,     295.8,   295.8,   295.8,
  295.4,     295.4,   295.4,   295.4,
  294.8,     294.8,   294.8,   294.8,
  294.6,     294.6,   294.6,   294.6,
  294.4,     294.4,   294.4,   294.4,
  293.85,    293.85,  293.85,  293.85,
  293.15,    293.15,  293.15,  293.15,
  292.55,    292.55,  292.55,  292.55,
  292.25,    292.25,  292.25,  292.25,
  292.1,     292.1,   292.1,   292.1,
  292.05,    292.05,  292.05,  292.05,
  292.2,     292.2,   292.2,   292.2,
  292.65,    292.65,  292.65,  292.65,
  293.35,    293.35,  293.35,  293.35,
  294.2,     294.2,   294.2,   294.2,
  295.1,     295.1,   295.1,   295.1,
  296,       296,     296,     296,
  296.95,    296.95,  296.95,  296.95,
  297.85,    297.85,  297.85,  297.85,
  298.65,    298.65,  298.65,  298.65,
  299.35,    299.35,  299.35,  299.35,
  300.05,    300.05,  300.05,  300.05,
  300.75,    300.75,  300.75,  300.75,
  301.25,    301.25,  301.25,  301.25,
  301.5,     301.5,   301.5,   301.5,
  301.8,     301.8,   301.8,   301.8,
  302.2,     302.2,   302.2,   302.2,
  302.5,     302.5,   302.5,   302.5,
  302.8,     302.8,   302.8,   302.8,
  303.1,     303.1,   303.1,   303.1,
  303.35,    303.35,  303.35,  303.35,
  303.45,    303.45,  303.45,  303.45,
  303.55,    303.55,  303.55,  303.55,
  303.65,    303.65,  303.65,  303.65,
  303.5,     303.5,   303.5,   303.5,
  303.2,     303.2,   303.2,   303.2,
  302.75,    302.75,  302.75,  302.75,
  302,       302,     302,     302,
  301,       301,     301,     301,
  299.9,     299.9,   299.9,   299.9,
  298.9,     298.9,   298.9,   298.9,
  298.1,     298.1,   298.1,   298.1,
  297.6,     297.6,   297.6,   297.6,
  297.3,     297.3,   297.3,   297.3,
  297,       297,     297,     297,
  296.65,    296.65,  296.65,  296.65,
  296.2,     296.2,   296.2,   296.2,
  295.75,    295.75,  295.75,  295.75,
  295.5,     295.5,   295.5,   295.5,
  295.5,     295.5,   295.5,   295.5,
  295.45,    295.45,  295.45,  295.45,
  295.2,     295.2,   295.2,   295.2,
  294.8,     294.8,   294.8,   294.8,
  294.25,    294.25,  294.25,  294.25,
  293.75,    293.75,  293.75,  293.75,
  293.5,     293.5,   293.5,   293.5,
  293.3,     293.3,   293.3,   293.3,
  292.8,     292.8,   292.8,   292.8,
  292.15,    292.15,  292.15,  292.15,
  291.9,     291.9,   291.9,   291.9,
  292.45,    292.45,  292.45,  292.45,
  293.75,    293.75,  293.75,  293.75,
  295.3,     295.3,   295.3,   295.3,
  296.75,    296.75,  296.75,  296.75,
  297.85,    297.85,  297.85,  297.85,
  298.7,     298.7,   298.7,   298.7,
  299.55,    299.55,  299.55,  299.55,
  300.35,    300.35,  300.35,  300.35,
  300.95,    300.95,  300.95,  300.95,
  301.45,    301.45,  301.45,  301.45,
  302.05,    302.05,  302.05,  302.05,
  302.4,     302.4,   302.4,   302.4,
  302.7,     302.7,   302.7,   302.7,
  302.9,     302.9,   302.9,   302.9,
  302.95,    302.95,  302.95,  302.95,
  303.1,     303.1,   303.1,   303.1,
  303.2,     303.2,   303.2,   303.2,
  303.35,    303.35,  303.35,  303.35,
  303.4,     303.4,   303.4,   303.4,
  303.25,    303.25,  303.25,  303.25,
  303,       303,     303,     303,
  302.65,    302.65,  302.65,  302.65,
  302.6,     302.6,   302.6,   302.6,
  302.7,     302.7,   302.7,   302.7,
  302.45,    302.45,  302.45,  302.45,
  302,       302,     302,     302,
  301.35,    301.35,  301.35,  301.35,
  300.25,    300.25,  300.25,  300.25,
  298.95,    298.95,  298.95,  298.95,
  298.05,    298.05,  298.05,  298.05,
  297.4,     297.4,   297.4,   297.4,
  296.65,    296.65,  296.65,  296.65,
  296.05,    296.05,  296.05,  296.05,
  295.65,    295.65,  295.65,  295.65,
  295.3,     295.3,   295.3,   295.3,
  295.15,    295.15,  295.15,  295.15,
  294.9,     294.9,   294.9,   294.9,
  294.4,     294.4,   294.4,   294.4,
  294.15,    294.15,  294.15,  294.15,
  293.95,    293.95,  293.95,  293.95,
  293.55,    293.55,  293.55,  293.55,
  293,       293,     293,     293,
  292.15,    292.15,  292.15,  292.15,
  291.35,    291.35,  291.35,  291.35,
  291.3,     291.3,   291.3,   291.3,
  291.6,     291.6,   291.6,   291.6,
  291.6,     291.6,   291.6,   291.6,
  291.5,     291.5,   291.5,   291.5,
  291.6,     291.6,   291.6,   291.6,
  292.6,     292.6,   292.6,   292.6,
  294.4,     294.4,   294.4,   294.4,
  296.15,    296.15,  296.15,  296.15,
  297.6,     297.6,   297.6,   297.6,
  298.85,    298.85,  298.85,  298.85,
  299.95,    299.95,  299.95,  299.95,
  300.9,     300.9,   300.9,   300.9,
  301.55,    301.55,  301.55,  301.55,
  302.3,     302.3,   302.3,   302.3,
  303.15,    303.15,  303.15,  303.15,
  303.65,    303.65,  303.65,  303.65,
  304.05,    304.05,  304.05,  304.05,
  304.2,     304.2,   304.2,   304.2,
  304.15,    304.15,  304.15,  304.15,
  304.2,     304.2,   304.2,   304.2,
  304.2,     304.2,   304.2,   304.2,
  304.15,    304.15,  304.15,  304.15,
  304,       304,     304,     304,
  303.9,     303.9,   303.9,   303.9,
  303.8,     303.8,   303.8,   303.8,
  303.55,    303.55,  303.55,  303.55,
  303.2,     303.2,   303.2,   303.2,
  302.65,    302.65,  302.65,  302.65,
  302.05,    302.05,  302.05,  302.05,
  301.35,    301.35,  301.35,  301.35,
  300.5,     300.5,   300.5,   300.5,
  299.1,     299.1,   299.1,   299.1,
  297.4,     297.4,   297.4,   297.4,
  296.2,     296.2,   296.2,   296.2,
  295.3,     295.3,   295.3,   295.3,
  294.5,     294.5,   294.5,   294.5,
  293.95,    293.95,  293.95,  293.95,
  293.5,     293.5,   293.5,   293.5,
  292.9,     292.9,   292.9,   292.9,
  292.3,     292.3,   292.3,   292.3,
  291.9,     291.9,   291.9,   291.9,
  291.35,    291.35,  291.35,  291.35,
  290.8,     290.8,   290.8,   290.8,
  290.55,    290.55,  290.55,  290.55,
  290.3,     290.3,   290.3,   290.3,
  289.9,     289.9,   289.9,   289.9,
  289.5,     289.5,   289.5,   289.5,
  289.3,     289.3,   289.3,   289.3,
  289.2,     289.2,   289.2,   289.2,
  289,       289,     289,     289,
  288.75,    288.75,  288.75,  288.75,
  288.75,    288.75,  288.75,  288.75,
  289.15,    289.15,  289.15,  289.15,
  289.5,     289.5,   289.5,   289.5,
  289.7,     289.7,   289.7,   289.7,
  290.05,    290.05,  290.05,  290.05,
  290.35,    290.35,  290.35,  290.35,
  290.6,     290.6,   290.6,   290.6,
  291.25,    291.25,  291.25,  291.25,
  292.6,     292.6,   292.6,   292.6,
  293.85,    293.85,  293.85,  293.85,
  294,       294,     294,     294,
  293.7,     293.7,   293.7,   293.7,
  293.6,     293.6,   293.6,   293.6,
  293.65,    293.65,  293.65,  293.65,
  294.05,    294.05,  294.05,  294.05,
  294.3,     294.3,   294.3,   294.3,
  294.3,     294.3,   294.3,   294.3,
  294.2,     294.2,   294.2,   294.2,
  293.85,    293.85,  293.85,  293.85,
  293.5,     293.5,   293.5,   293.5,
  293.45,    293.45,  293.45,  293.45,
  293.85,    293.85,  293.85,  293.85,
  294.4,     294.4,   294.4,   294.4,
  294.45,    294.45,  294.45,  294.45,
  294,       294,     294,     294,
  293.55,    293.55,  293.55,  293.55,
  293.05,    293.05,  293.05,  293.05,
  292.75,    292.75,  292.75,  292.75,
  292.65,    292.65,  292.65,  292.65,
  292.5,     292.5,   292.5,   292.5,
  292.35,    292.35,  292.35,  292.35,
  292.1,     292.1,   292.1,   292.1,
  291.85,    291.85,  291.85,  291.85,
  291.7,     291.7,   291.7,   291.7,
  291.5,     291.5,   291.5,   291.5,
  291.2,     291.2,   291.2,   291.2,
  291,       291,     291,     291,
  290.7,     290.7,   290.7,   290.7,
  290.3,     290.3,   290.3,   290.3,
  289.95,    289.95,  289.95,  289.95,
  289.45,    289.45,  289.45,  289.45,
  288.95,    288.95,  288.95,  288.95,
  288.7,     288.7,   288.7,   288.7,
  288.5,     288.5,   288.5,   288.5,
  288.25,    288.25,  288.25,  288.25,
  288.05,    288.05,  288.05,  288.05,
  288,       288,     288,     288,
  288.1,     288.1,   288.1,   288.1,
  288.25,    288.25,  288.25,  288.25,
  288.45,    288.45,  288.45,  288.45,
  288.85,    288.85,  288.85,  288.85,
  289.7,     289.7,   289.7,   289.7,
  290.9,     290.9,   290.9,   290.9,
  291.8,     291.8,   291.8,   291.8,
  292.3,     292.3,   292.3,   292.3,
  292.8,     292.8,   292.8,   292.8,
  293.4,     293.4,   293.4,   293.4,
  294,       294,     294,     294,
  294.5,     294.5,   294.5,   294.5,
  295,       295,     295,     295,
  295.5,     295.5,   295.5,   295.5,
  295.9,     295.9,   295.9,   295.9,
  296.4,     296.4,   296.4,   296.4,
  296.75,    296.75,  296.75,  296.75,
  296.7,     296.7,   296.7,   296.7,
  296.75,    296.75,  296.75,  296.75,
  297,       297,     297,     297,
  297.15,    297.15,  297.15,  297.15,
  297.3,     297.3,   297.3,   297.3,
  297.15,    297.15,  297.15,  297.15,
  296.6,     296.6,   296.6,   296.6,
  296.25,    296.25,  296.25,  296.25,
  295.9,     295.9,   295.9,   295.9,
  295.35,    295.35,  295.35,  295.35,
  294.65,    294.65,  294.65,  294.65,
  293.8,     293.8,   293.8,   293.8,
  292.95,    292.95,  292.95,  292.95,
  292.2,     292.2,   292.2,   292.2,
  291.6,     291.6,   291.6,   291.6,
  291.05,    291.05,  291.05,  291.05,
  290.5,     290.5,   290.5,   290.5,
  290.05,    290.05,  290.05,  290.05,
  289.7,     289.7,   289.7,   289.7,
  289.45,    289.45,  289.45,  289.45,
  289.1,     289.1,   289.1,   289.1,
  288.9,     288.9,   288.9,   288.9,
  288.75,    288.75,  288.75,  288.75,
  288.1,     288.1,   288.1,   288.1,
  287.2,     287.2,   287.2,   287.2,
  286.35,    286.35,  286.35,  286.35,
  286.55,    286.55,  286.55,  286.55,
  286.9,     286.9,   286.9,   286.9,
  286.05,    286.05,  286.05,  286.05,
  285.75,    285.75,  285.75,  285.75,
  286.15,    286.15,  286.15,  286.15,
  286.05,    286.05,  286.05,  286.05,
  286.35,    286.35,  286.35,  286.35,
  286.75,    286.75,  286.75,  286.75,
  286.8,     286.8,   286.8,   286.8,
  287.95,    287.95,  287.95,  287.95,
  289.75,    289.75,  289.75,  289.75,
  290.8,     290.8,   290.8,   290.8,
  291.75,    291.75,  291.75,  291.75,
  293.1,     293.1,   293.1,   293.1,
  294.15,    294.15,  294.15,  294.15,
  294.85,    294.85,  294.85,  294.85,
  295.1,     295.1,   295.1,   295.1,
  295.25,    295.25,  295.25,  295.25,
  295.95,    295.95,  295.95,  295.95,
  296.65,    296.65,  296.65,  296.65,
  296.75,    296.75,  296.75,  296.75,
  296.65,    296.65,  296.65,  296.65,
  296.75,    296.75,  296.75,  296.75,
  297.15,    297.15,  297.15,  297.15,
  297.25,    297.25,  297.25,  297.25,
  297.4,     297.4,   297.4,   297.4,
  297.5,     297.5,   297.5,   297.5,
  297.5,     297.5,   297.5,   297.5,
  297.7,     297.7,   297.7,   297.7,
  297.35,    297.35,  297.35,  297.35,
  296.8,     296.8,   296.8,   296.8,
  296.35,    296.35,  296.35,  296.35,
  295.95,    295.95,  295.95,  295.95,
  295.45,    295.45,  295.45,  295.45,
  294.75,    294.75,  294.75,  294.75,
  293.85,    293.85,  293.85,  293.85,
  293.1,     293.1,   293.1,   293.1,
  292.55,    292.55,  292.55,  292.55,
  292.15,    292.15,  292.15,  292.15,
  292.05,    292.05,  292.05,  292.05,
  291.9,     291.9,   291.9,   291.9,
  291.6,     291.6,   291.6,   291.6,
  291.2,     291.2,   291.2,   291.2,
  290.9,     290.9,   290.9,   290.9,
  290.6,     290.6,   290.6,   290.6,
  290.15,    290.15,  290.15,  290.15,
  289.95,    289.95,  289.95,  289.95,
  289.8,     289.8,   289.8,   289.8,
  289.45,    289.45,  289.45,  289.45,
  289.2,     289.2,   289.2,   289.2,
  288.9,     288.9,   288.9,   288.9,
  288.55,    288.55,  288.55,  288.55,
  288.25,    288.25,  288.25,  288.25,
  288,       288,     288,     288,
  287.9,     287.9,   287.9,   287.9,
  288.15,    288.15,  288.15,  288.15,
  288.9,     288.9,   288.9,   288.9,
  289.95,    289.95,  289.95,  289.95,
  291.5,     291.5,   291.5,   291.5,
  293.3,     293.3,   293.3,   293.3,
  295,       295,     295,     295,
  296.3,     296.3,   296.3,   296.3,
  297.1,     297.1,   297.1,   297.1,
  297.75,    297.75,  297.75,  297.75,
  298.4,     298.4,   298.4,   298.4,
  299.15,    299.15,  299.15,  299.15,
  299.65,    299.65,  299.65,  299.65,
  299.8,     299.8,   299.8,   299.8,
  300.2,     300.2,   300.2,   300.2,
  300.6,     300.6,   300.6,   300.6,
  300.75,    300.75,  300.75,  300.75,
  300.9,     300.9,   300.9,   300.9,
  301.05,    301.05,  301.05,  301.05,
  301.2,     301.2,   301.2,   301.2,
  301.15,    301.15,  301.15,  301.15,
  300.7,     300.7,   300.7,   300.7,
  300.25,    300.25,  300.25,  300.25,
  299.6,     299.6,   299.6,   299.6,
  298.8,     298.8,   298.8,   298.8,
  298.55,    298.55,  298.55,  298.55,
  298.3,     298.3,   298.3,   298.3,
  297.65,    297.65,  297.65,  297.65,
  296.75,    296.75,  296.75,  296.75,
  295.8,     295.8,   295.8,   295.8,
  295.05,    295.05,  295.05,  295.05,
  294.4,     294.4,   294.4,   294.4,
  294,       294,     294,     294,
  293.9,     293.9,   293.9,   293.9,
  293.75,    293.75,  293.75,  293.75,
  293.35,    293.35,  293.35,  293.35,
  292.75,    292.75,  292.75,  292.75,
  292.45,    292.45,  292.45,  292.45,
  291.6,     291.6,   291.6,   291.6,
  290.75,    290.75,  290.75,  290.75,
  290.65,    290.65,  290.65,  290.65,
  290.6,     290.6,   290.6,   290.6,
  290.4,     290.4,   290.4,   290.4,
  289.9,     289.9,   289.9,   289.9,
  289.75,    289.75,  289.75,  289.75,
  289.9,     289.9,   289.9,   289.9,
  289.8,     289.8,   289.8,   289.8,
  289.5,     289.5,   289.5,   289.5,
  289.6,     289.6,   289.6,   289.6,
  290,       290,     290,     290,
  290.4,     290.4,   290.4,   290.4,
  291.45,    291.45,  291.45,  291.45,
  293.15,    293.15,  293.15,  293.15,
  294.8,     294.8,   294.8,   294.8,
  296.35,    296.35,  296.35,  296.35,
  297.6,     297.6,   297.6,   297.6,
  298.25,    298.25,  298.25,  298.25,
  298.85,    298.85,  298.85,  298.85,
  299.45,    299.45,  299.45,  299.45,
  299.75,    299.75,  299.75,  299.75,
  299.95,    299.95,  299.95,  299.95,
  300.15,    300.15,  300.15,  300.15,
  300.5,     300.5,   300.5,   300.5,
  301,       301,     301,     301,
  301.3,     301.3,   301.3,   301.3,
  301.2,     301.2,   301.2,   301.2,
  301.2,     301.2,   301.2,   301.2,
  301.4,     301.4,   301.4,   301.4,
  301.45,    301.45,  301.45,  301.45,
  301.35,    301.35,  301.35,  301.35,
  301.1,     301.1,   301.1,   301.1,
  300.95,    300.95,  300.95,  300.95,
  300.8,     300.8,   300.8,   300.8,
  300.4,     300.4,   300.4,   300.4,
  299.8,     299.8,   299.8,   299.8,
  299.2,     299.2,   299.2,   299.2,
  298.6,     298.6,   298.6,   298.6,
  297.8,     297.8,   297.8,   297.8,
  296.8,     296.8,   296.8,   296.8,
  295.65,    295.65,  295.65,  295.65,
  294.6,     294.6,   294.6,   294.6,
  294,       294,     294,     294,
  293.55,    293.55,  293.55,  293.55,
  293.1,     293.1,   293.1,   293.1,
  292.75,    292.75,  292.75,  292.75,
  292.4,     292.4,   292.4,   292.4,
  292.15,    292.15,  292.15,  292.15,
  291.9,     291.9,   291.9,   291.9,
  291.6,     291.6,   291.6,   291.6,
  291.35,    291.35,  291.35,  291.35,
  291.15,    291.15,  291.15,  291.15,
  290.8,     290.8,   290.8,   290.8,
  290.35,    290.35,  290.35,  290.35,
  289.8,     289.8,   289.8,   289.8,
  289.45,    289.45,  289.45,  289.45,
  289.3,     289.3,   289.3,   289.3,
  289.05,    289.05,  289.05,  289.05,
  289.2,     289.2,   289.2,   289.2,
  290,       290,     290,     290,
  291.4,     291.4,   291.4,   291.4,
  292.95,    292.95,  292.95,  292.95,
  293.85,    293.85,  293.85,  293.85,
  294.9,     294.9,   294.9,   294.9,
  296.2,     296.2,   296.2,   296.2,
  296.7,     296.7,   296.7,   296.7,
  297.05,    297.05,  297.05,  297.05,
  297.5,     297.5,   297.5,   297.5,
  298,       298,     298,     298,
  298.3,     298.3,   298.3,   298.3,
  298.4,     298.4,   298.4,   298.4,
  298.75,    298.75,  298.75,  298.75,
  299,       299,     299,     299,
  299.05,    299.05,  299.05,  299.05,
  298.9,     298.9,   298.9,   298.9,
  298.7,     298.7,   298.7,   298.7,
  298.55,    298.55,  298.55,  298.55,
  298.35,    298.35,  298.35,  298.35,
  298.15,    298.15,  298.15,  298.15,
  297.85,    297.85,  297.85,  297.85,
  297.5,     297.5,   297.5,   297.5,
  296.85,    296.85,  296.85,  296.85,
  295.95,    295.95,  295.95,  295.95,
  295.1,     295.1,   295.1,   295.1,
  294.2,     294.2,   294.2,   294.2,
  293.45,    293.45,  293.45,  293.45,
  292.85,    292.85,  292.85,  292.85,
  292.25,    292.25,  292.25,  292.25,
  291.65,    291.65,  291.65,  291.65,
  291.05,    291.05,  291.05,  291.05,
  290.55,    290.55,  290.55,  290.55,
  290.2,     290.2,   290.2,   290.2,
  289.8,     289.8,   289.8,   289.8,
  289.4,     289.4,   289.4,   289.4,
  289.05,    289.05,  289.05,  289.05,
  288.65,    288.65,  288.65,  288.65,
  288.45,    288.45,  288.45,  288.45,
  288.4,     288.4,   288.4,   288.4,
  288.55,    288.55,  288.55,  288.55,
  288.9,     288.9,   288.9,   288.9,
  288.9,     288.9,   288.9,   288.9,
  288.6,     288.6,   288.6,   288.6,
  288.55,    288.55,  288.55,  288.55,
  288.7,     288.7,   288.7,   288.7,
  288.65,    288.65,  288.65,  288.65,
  288.55,    288.55,  288.55,  288.55,
  288.7,     288.7,   288.7,   288.7,
  289.3,     289.3,   289.3,   289.3,
  290.45,    290.45,  290.45,  290.45,
  291.8,     291.8,   291.8,   291.8,
  293.1,     293.1,   293.1,   293.1,
  294.4,     294.4,   294.4,   294.4,
  295.55,    295.55,  295.55,  295.55,
  296.05,    296.05,  296.05,  296.05,
  295.95,    295.95,  295.95,  295.95,
  296,       296,     296,     296,
  296.4,     296.4,   296.4,   296.4,
  296.65,    296.65,  296.65,  296.65,
  296.65,    296.65,  296.65,  296.65,
  296.8,     296.8,   296.8,   296.8,
  297.15,    297.15,  297.15,  297.15,
  297.6,     297.6,   297.6,   297.6,
  298,       298,     298,     298,
  298.15,    298.15,  298.15,  298.15,
  298.35,    298.35,  298.35,  298.35,
  298.55,    298.55,  298.55,  298.55,
  298.5,     298.5,   298.5,   298.5,
  298.35,    298.35,  298.35,  298.35,
  298.15,    298.15,  298.15,  298.15,
  298.05,    298.05,  298.05,  298.05,
  297.9,     297.9,   297.9,   297.9,
  297.55,    297.55,  297.55,  297.55,
  297.15,    297.15,  297.15,  297.15,
  296.5,     296.5,   296.5,   296.5,
  295.75,    295.75,  295.75,  295.75,
  295,       295,     295,     295,
  293.9,     293.9,   293.9,   293.9,
  293.05,    293.05,  293.05,  293.05,
  292.65,    292.65,  292.65,  292.65,
  291.85,    291.85,  291.85,  291.85,
  291.4,     291.4,   291.4,   291.4,
  291.5,     291.5,   291.5,   291.5,
  291.6,     291.6,   291.6,   291.6,
  291,       291,     291,     291,
  290.25,    290.25,  290.25,  290.25,
  290.45,    290.45,  290.45,  290.45,
  290.7,     290.7,   290.7,   290.7,
  290.45,    290.45,  290.45,  290.45,
  289.9,     289.9,   289.9,   289.9,
  289.7,     289.7,   289.7,   289.7,
  289.7,     289.7,   289.7,   289.7,
  289.45,    289.45,  289.45,  289.45,
  289.35,    289.35,  289.35,  289.35,
  289.6,     289.6,   289.6,   289.6,
  289.95,    289.95,  289.95,  289.95,
  290.25,    290.25,  290.25,  290.25,
  290.8,     290.8,   290.8,   290.8,
  291.85,    291.85,  291.85,  291.85,
  293.15,    293.15,  293.15,  293.15,
  294.4,     294.4,   294.4,   294.4,
  295.4,     295.4,   295.4,   295.4,
  296.35,    296.35,  296.35,  296.35,
  297.15,    297.15,  297.15,  297.15,
  297.7,     297.7,   297.7,   297.7,
  298.2,     298.2,   298.2,   298.2,
  298.65,    298.65,  298.65,  298.65,
  299,       299,     299,     299,
  299.1,     299.1,   299.1,   299.1,
  299.3,     299.3,   299.3,   299.3,
  299.7,     299.7,   299.7,   299.7,
  300.05,    300.05,  300.05,  300.05,
  300.3,     300.3,   300.3,   300.3,
  300.3,     300.3,   300.3,   300.3,
  300.3,     300.3,   300.3,   300.3,
  300.35,    300.35,  300.35,  300.35,
  300.3,     300.3,   300.3,   300.3,
  300.25,    300.25,  300.25,  300.25,
  300.2,     300.2,   300.2,   300.2,
  299.9,     299.9,   299.9,   299.9,
  299.3,     299.3,   299.3,   299.3,
  298.75,    298.75,  298.75,  298.75,
  298.3,     298.3,   298.3,   298.3,
  297.75,    297.75,  297.75,  297.75,
  296.5,     296.5,   296.5,   296.5,
  295.5,     295.5,   295.5,   295.5,
  295.2,     295.2,   295.2,   295.2,
  294.6,     294.6,   294.6,   294.6,
  294.15,    294.15,  294.15,  294.15,
  294,       294,     294,     294,
  294,       294,     294,     294,
  294,       294,     294,     294,
  293.8,     293.8,   293.8,   293.8,
  293.6,     293.6,   293.6,   293.6,
  293.4,     293.4,   293.4,   293.4,
  293.35,    293.35,  293.35,  293.35,
  293.5,     293.5,   293.5,   293.5,
  293.55,    293.55,  293.55,  293.55,
  293.5,     293.5,   293.5,   293.5,
  293.2,     293.2,   293.2,   293.2,
  292.7,     292.7,   292.7,   292.7,
  292.4,     292.4,   292.4,   292.4,
  292.3,     292.3,   292.3,   292.3,
  292.3,     292.3,   292.3,   292.3,
  292.5,     292.5,   292.5,   292.5,
  292.95,    292.95,  292.95,  292.95,
  293.4,     293.4,   293.4,   293.4,
  293.65,    293.65,  293.65,  293.65,
  293.65,    293.65,  293.65,  293.65,
  293.45,    293.45,  293.45,  293.45,
  293.05,    293.05,  293.05,  293.05,
  292.7,     292.7,   292.7,   292.7,
  292.25,    292.25,  292.25,  292.25,
  291.95,    291.95,  291.95,  291.95,
  292.2,     292.2,   292.2,   292.2,
  292.35,    292.35,  292.35,  292.35,
  292.3,     292.3,   292.3,   292.3,
  292.2,     292.2,   292.2,   292.2,
  292.15,    292.15,  292.15,  292.15,
  292.15,    292.15,  292.15,  292.15,
  292.15,    292.15,  292.15,  292.15,
  292.25,    292.25,  292.25,  292.25,
  292.45,    292.45,  292.45,  292.45,
  292.6,     292.6,   292.6,   292.6,
  292.7,     292.7,   292.7,   292.7,
  292.8,     292.8,   292.8,   292.8,
  292.9,     292.9,   292.9,   292.9,
  292.95,    292.95,  292.95,  292.95,
  292.95,    292.95,  292.95,  292.95,
  292.95,    292.95,  292.95,  292.95,
  292.9,     292.9,   292.9,   292.9,
  292.8,     292.8,   292.8,   292.8,
  292.7,     292.7,   292.7,   292.7,
  292.65,    292.65,  292.65,  292.65,
  292.6,     292.6,   292.6,   292.6,
  292.5,     292.5,   292.5,   292.5,
  292.45,    292.45,  292.45,  292.45,
  292.45,    292.45,  292.45,  292.45,
  292.45,    292.45,  292.45,  292.45,
  292.45,    292.45,  292.45,  292.45,
  292.4,     292.4,   292.4,   292.4,
  292.3,     292.3,   292.3,   292.3,
  292.2,     292.2,   292.2,   292.2,
  292.15,    292.15,  292.15,  292.15,
  292.1,     292.1,   292.1,   292.1,
  292.05,    292.05,  292.05,  292.05,
  292.05,    292.05,  292.05,  292.05,
  292.05,    292.05,  292.05,  292.05,
  292.05,    292.05,  292.05,  292.05,
  292,       292,     292,     292,
  291.95,    291.95,  291.95,  291.95,
  291.9,     291.9,   291.9,   291.9,
  291.85,    291.85,  291.85,  291.85,
  291.8,     291.8,   291.8,   291.8,
  291.7,     291.7,   291.7,   291.7,
  291.8,     291.8,   291.8,   291.8,
  292.1,     292.1,   292.1,   292.1,
  292.4,     292.4,   292.4,   292.4,
  292.85,    292.85,  292.85,  292.85,
  293.35,    293.35,  293.35,  293.35,
  293.85,    293.85,  293.85,  293.85,
  294.45,    294.45,  294.45,  294.45,
  295,       295,     295,     295,
  295.45,    295.45,  295.45,  295.45,
  295.9,     295.9,   295.9,   295.9,
  296.3,     296.3,   296.3,   296.3,
  296.55,    296.55,  296.55,  296.55,
  296.75,    296.75,  296.75,  296.75,
  296.95,    296.95,  296.95,  296.95,
  297.15,    297.15,  297.15,  297.15,
  297.4,     297.4,   297.4,   297.4,
  297.6,     297.6,   297.6,   297.6,
  297.6,     297.6,   297.6,   297.6,
  297.4,     297.4,   297.4,   297.4,
  297.1,     297.1,   297.1,   297.1,
  296.95,    296.95,  296.95,  296.95,
  296.9,     296.9,   296.9,   296.9,
  296.7,     296.7,   296.7,   296.7,
  296.25,    296.25,  296.25,  296.25,
  295.6,     295.6,   295.6,   295.6,
  295.2,     295.2,   295.2,   295.2,
  294.95,    294.95,  294.95,  294.95,
  294.6,     294.6,   294.6,   294.6,
  294.4,     294.4,   294.4,   294.4,
  294.25,    294.25,  294.25,  294.25,
  294.25,    294.25,  294.25,  294.25,
  294.45,    294.45,  294.45,  294.45,
  294.6,     294.6,   294.6,   294.6,
  294.65,    294.65,  294.65,  294.65,
  294.6,     294.6,   294.6,   294.6,
  294.45,    294.45,  294.45,  294.45,
  294.25,    294.25,  294.25,  294.25,
  294.1,     294.1,   294.1,   294.1,
  293.95,    293.95,  293.95,  293.95,
  293.85,    293.85,  293.85,  293.85,
  293.85,    293.85,  293.85,  293.85,
  293.75,    293.75,  293.75,  293.75,
  293.55,    293.55,  293.55,  293.55,
  293.4,     293.4,   293.4,   293.4,
  293.5,     293.5,   293.5,   293.5,
  294.05,    294.05,  294.05,  294.05,
  294.85,    294.85,  294.85,  294.85,
  295.35,    295.35,  295.35,  295.35,
  295.75,    295.75,  295.75,  295.75,
  296.25,    296.25,  296.25,  296.25,
  296.65,    296.65,  296.65,  296.65,
  297,       297,     297,     297,
  297.35,    297.35,  297.35,  297.35,
  297.9,     297.9,   297.9,   297.9,
  298.55,    298.55,  298.55,  298.55,
  299.15,    299.15,  299.15,  299.15,
  299.65,    299.65,  299.65,  299.65,
  300.05,    300.05,  300.05,  300.05,
  300.4,     300.4,   300.4,   300.4,
  300.65,    300.65,  300.65,  300.65,
  300.75,    300.75,  300.75,  300.75,
  300.8,     300.8,   300.8,   300.8,
  300.85,    300.85,  300.85,  300.85,
  300.8,     300.8,   300.8,   300.8,
  300.75,    300.75,  300.75,  300.75,
  300.65,    300.65,  300.65,  300.65,
  300.35,    300.35,  300.35,  300.35,
  300.05,    300.05,  300.05,  300.05,
  299.8,     299.8,   299.8,   299.8,
  299.3,     299.3,   299.3,   299.3,
  298.8,     298.8,   298.8,   298.8,
  298.4,     298.4,   298.4,   298.4,
  297.4,     297.4,   297.4,   297.4,
  296.05,    296.05,  296.05,  296.05,
  295.4,     295.4,   295.4,   295.4,
  295.25,    295.25,  295.25,  295.25,
  295.1,     295.1,   295.1,   295.1,
  295.1,     295.1,   295.1,   295.1,
  295.3,     295.3,   295.3,   295.3,
  295.5,     295.5,   295.5,   295.5,
  295.15,    295.15,  295.15,  295.15,
  293.6,     293.6,   293.6,   293.6,
  292.4,     292.4,   292.4,   292.4,
  292.45,    292.45,  292.45,  292.45,
  292.65,    292.65,  292.65,  292.65,
  292.8,     292.8,   292.8,   292.8,
  292.85,    292.85,  292.85,  292.85,
  292.8,     292.8,   292.8,   292.8,
  292.6,     292.6,   292.6,   292.6,
  292.35,    292.35,  292.35,  292.35,
  292.2,     292.2,   292.2,   292.2,
  292.15,    292.15,  292.15,  292.15,
  292.25,    292.25,  292.25,  292.25,
  292.5,     292.5,   292.5,   292.5,
  292.9,     292.9,   292.9,   292.9,
  293.45,    293.45,  293.45,  293.45,
  294.1,     294.1,   294.1,   294.1,
  294.75,    294.75,  294.75,  294.75,
  295.25,    295.25,  295.25,  295.25,
  295.95,    295.95,  295.95,  295.95,
  296.9,     296.9,   296.9,   296.9,
  297.55,    297.55,  297.55,  297.55,
  298.15,    298.15,  298.15,  298.15,
  298.95,    298.95,  298.95,  298.95,
  299.75,    299.75,  299.75,  299.75,
  300.8,     300.8,   300.8,   300.8,
  301.8,     301.8,   301.8,   301.8,
  302.6,     302.6,   302.6,   302.6,
  303.25,    303.25,  303.25,  303.25,
  303.55,    303.55,  303.55,  303.55,
  303.3,     303.3,   303.3,   303.3,
  302.65,    302.65,  302.65,  302.65,
  298.6,     298.6,   298.6,   298.6,
  293.65,    293.65,  293.65,  293.65,
  292.45,    292.45,  292.45,  292.45,
  292.45,    292.45,  292.45,  292.45,
  292.55,    292.55,  292.55,  292.55,
  292.65,    292.65,  292.65,  292.65,
  292.65,    292.65,  292.65,  292.65,
  292.65,    292.65,  292.65,  292.65,
  292.65,    292.65,  292.65,  292.65,
  292.6,     292.6,   292.6,   292.6,
  292.5,     292.5,   292.5,   292.5,
  292.45,    292.45,  292.45,  292.45,
  292.25,    292.25,  292.25,  292.25,
  291.9,     291.9,   291.9,   291.9,
  291.6,     291.6,   291.6,   291.6,
  291.35,    291.35,  291.35,  291.35,
  291.25,    291.25,  291.25,  291.25,
  291.25,    291.25,  291.25,  291.25,
  291.2,     291.2,   291.2,   291.2,
  291.15,    291.15,  291.15,  291.15,
  291.1,     291.1,   291.1,   291.1,
  290.95,    290.95,  290.95,  290.95,
  290.8,     290.8,   290.8,   290.8,
  290.75,    290.75,  290.75,  290.75,
  290.85,    290.85,  290.85,  290.85,
  291,       291,     291,     291,
  291.1,     291.1,   291.1,   291.1,
  291.15,    291.15,  291.15,  291.15,
  291.15,    291.15,  291.15,  291.15,
  291.15,    291.15,  291.15,  291.15,
  291.15,    291.15,  291.15,  291.15,
  291.25,    291.25,  291.25,  291.25,
  291.5,     291.5,   291.5,   291.5,
  291.8,     291.8,   291.8,   291.8,
  292.1,     292.1,   292.1,   292.1,
  292.4,     292.4,   292.4,   292.4,
  292.7,     292.7,   292.7,   292.7,
  293.05,    293.05,  293.05,  293.05,
  293.35,    293.35,  293.35,  293.35,
  293.4,     293.4,   293.4,   293.4,
  293.35,    293.35,  293.35,  293.35,
  293.7,     293.7,   293.7,   293.7,
  294.05,    294.05,  294.05,  294.05,
  294,       294,     294,     294,
  293.9,     293.9,   293.9,   293.9,
  293.8,     293.8,   293.8,   293.8,
  293.7,     293.7,   293.7,   293.7,
  293.45,    293.45,  293.45,  293.45,
  293.2,     293.2,   293.2,   293.2,
  293.15,    293.15,  293.15,  293.15,
  293.15,    293.15,  293.15,  293.15,
  293.15,    293.15,  293.15,  293.15,
  293.15,    293.15,  293.15,  293.15,
  292.9,     292.9,   292.9,   292.9,
  292.4,     292.4,   292.4,   292.4,
  291.8,     291.8,   291.8,   291.8,
  291.2,     291.2,   291.2,   291.2,
  290.85,    290.85,  290.85,  290.85,
  290.6,     290.6,   290.6,   290.6,
  290.3,     290.3,   290.3,   290.3,
  290.05,    290.05,  290.05,  290.05,
  289.95,    289.95,  289.95,  289.95,
  289.9,     289.9,   289.9,   289.9,
  289.55,    289.55,  289.55,  289.55,
  288.7,     288.7,   288.7,   288.7,
  288.2,     288.2,   288.2,   288.2,
  288.35,    288.35,  288.35,  288.35,
  288.45,    288.45,  288.45,  288.45,
  288.5,     288.5,   288.5,   288.5,
  288.5,     288.5,   288.5,   288.5,
  288.45,    288.45,  288.45,  288.45,
  288.5,     288.5,   288.5,   288.5,
  288.35,    288.35,  288.35,  288.35,
  288.05,    288.05,  288.05,  288.05,
  288.05,    288.05,  288.05,  288.05,
  288.35,    288.35,  288.35,  288.35,
  288.7,     288.7,   288.7,   288.7,
  288.95,    288.95,  288.95,  288.95,
  289.25,    289.25,  289.25,  289.25,
  289.55,    289.55,  289.55,  289.55,
  289.85,    289.85,  289.85,  289.85,
  290.3,     290.3,   290.3,   290.3,
  290.6,     290.6,   290.6,   290.6,
  291.15,    291.15,  291.15,  291.15,
  292.45,    292.45,  292.45,  292.45,
  293.7,     293.7,   293.7,   293.7,
  294.45,    294.45,  294.45,  294.45,
  295.05,    295.05,  295.05,  295.05,
  295.6,     295.6,   295.6,   295.6,
  296.15,    296.15,  296.15,  296.15,
  296.5,     296.5,   296.5,   296.5,
  296.75,    296.75,  296.75,  296.75,
  297,       297,     297,     297,
  297.15,    297.15,  297.15,  297.15,
  297.05,    297.05,  297.05,  297.05,
  296.65,    296.65,  296.65,  296.65,
  294.5,     294.5,   294.5,   294.5,
  291.95,    291.95,  291.95,  291.95,
  291.2,     291.2,   291.2,   291.2,
  291.1,     291.1,   291.1,   291.1,
  291.25,    291.25,  291.25,  291.25,
  291.3,     291.3,   291.3,   291.3,
  291.1,     291.1,   291.1,   291.1,
  290.9,     290.9,   290.9,   290.9,
  290.75,    290.75,  290.75,  290.75,
  290.5,     290.5,   290.5,   290.5,
  290.4,     290.4,   290.4,   290.4,
  290.5,     290.5,   290.5,   290.5,
  290.65,    290.65,  290.65,  290.65,
  290.8,     290.8,   290.8,   290.8,
  290.95,    290.95,  290.95,  290.95,
  291.05,    291.05,  291.05,  291.05,
  291.05,    291.05,  291.05,  291.05,
  291,       291,     291,     291,
  290.85,    290.85,  290.85,  290.85,
  290.65,    290.65,  290.65,  290.65,
  290.5,     290.5,   290.5,   290.5,
  290.35,    290.35,  290.35,  290.35,
  290.2,     290.2,   290.2,   290.2,
  290.1,     290.1,   290.1,   290.1,
  290,       290,     290,     290,
  289.9,     289.9,   289.9,   289.9,
  289.85,    289.85,  289.85,  289.85,
  289.75,    289.75,  289.75,  289.75,
  289.65,    289.65,  289.65,  289.65,
  289.65,    289.65,  289.65,  289.65,
  289.65,    289.65,  289.65,  289.65,
  289.7,     289.7,   289.7,   289.7,
  289.8,     289.8,   289.8,   289.8,
  289.9,     289.9,   289.9,   289.9,
  289.9,     289.9,   289.9,   289.9,
  289.9,     289.9,   289.9,   289.9,
  289.75,    289.75,  289.75,  289.75,
  289.4,     289.4,   289.4,   289.4,
  289.35,    289.35,  289.35,  289.35,
  289.65,    289.65,  289.65,  289.65,
  290.05,    290.05,  290.05,  290.05,
  290.25,    290.25,  290.25,  290.25,
  290.25,    290.25,  290.25,  290.25,
  290.25,    290.25,  290.25,  290.25,
  290.1,     290.1,   290.1,   290.1,
  290.15,    290.15,  290.15,  290.15,
  290.3,     290.3,   290.3,   290.3,
  290.3,     290.3,   290.3,   290.3,
  290.6,     290.6,   290.6,   290.6,
  290.9,     290.9,   290.9,   290.9,
  290.75,    290.75,  290.75,  290.75,
  290.4,     290.4,   290.4,   290.4,
  290.2,     290.2,   290.2,   290.2,
  290.15,    290.15,  290.15,  290.15,
  289.8,     289.8,   289.8,   289.8,
  289,       289,     289,     289,
  288.25,    288.25,  288.25,  288.25,
  287.8,     287.8,   287.8,   287.8,
  287.6,     287.6,   287.6,   287.6,
  287.5,     287.5,   287.5,   287.5,
  287.5,     287.5,   287.5,   287.5,
  287.85,    287.85,  287.85,  287.85,
  288.15,    288.15,  288.15,  288.15,
  288.1,     288.1,   288.1,   288.1,
  288.1,     288.1,   288.1,   288.1,
  288.05,    288.05,  288.05,  288.05,
  287.85,    287.85,  287.85,  287.85,
  287.75,    287.75,  287.75,  287.75,
  287.85,    287.85,  287.85,  287.85,
  287.95,    287.95,  287.95,  287.95,
  287.85,    287.85,  287.85,  287.85,
  287.75,    287.75,  287.75,  287.75,
  287.75,    287.75,  287.75,  287.75,
  287.7,     287.7,   287.7,   287.7,
  287.75,    287.75,  287.75,  287.75,
  287.85,    287.85,  287.85,  287.85,
  287.9,     287.9,   287.9,   287.9,
  288,       288,     288,     288,
  288.2,     288.2,   288.2,   288.2,
  288.55,    288.55,  288.55,  288.55,
  288.9,     288.9,   288.9,   288.9,
  289.1,     289.1,   289.1,   289.1,
  289.3,     289.3,   289.3,   289.3,
  289.6,     289.6,   289.6,   289.6,
  290,       290,     290,     290,
  290.3,     290.3,   290.3,   290.3,
  290.6,     290.6,   290.6,   290.6,
  290.85,    290.85,  290.85,  290.85,
  290.75,    290.75,  290.75,  290.75,
  290.15,    290.15,  290.15,  290.15,
  290.15,    290.15,  290.15,  290.15,
  290.35,    290.35,  290.35,  290.35,
  290.4,     290.4,   290.4,   290.4,
  289.8,     289.8,   289.8,   289.8,
  289.25,    289.25,  289.25,  289.25,
  290.3,     290.3,   290.3,   290.3,
  290.75,    290.75,  290.75,  290.75,
  290.3,     290.3,   290.3,   290.3,
  289.85,    289.85,  289.85,  289.85,
  289,       289,     289,     289,
  288.1,     288.1,   288.1,   288.1,
  287.75,    287.75,  287.75,  287.75,
  287.35,    287.35,  287.35,  287.35,
  286.9,     286.9,   286.9,   286.9,
  286.85,    286.85,  286.85,  286.85,
  286.6,     286.6,   286.6,   286.6,
  286.05,    286.05,  286.05,  286.05,
  285.7,     285.7,   285.7,   285.7,
  285.45,    285.45,  285.45,  285.45,
  285.4,     285.4,   285.4,   285.4,
  285.45,    285.45,  285.45,  285.45,
  285.4,     285.4,   285.4,   285.4,
  285.15,    285.15,  285.15,  285.15,
  284.85,    284.85,  284.85,  284.85,
  284.35,    284.35,  284.35,  284.35,
  283.8,     283.8,   283.8,   283.8,
  283.6,     283.6,   283.6,   283.6,
  283.45,    283.45,  283.45,  283.45,
  283.35,    283.35,  283.35,  283.35,
  283.4,     283.4,   283.4,   283.4,
  283.55,    283.55,  283.55,  283.55,
  283.75,    283.75,  283.75,  283.75,
  283.9,     283.9,   283.9,   283.9,
  284,       284,     284,     284,
  284.3,     284.3,   284.3,   284.3,
  284.85,    284.85,  284.85,  284.85,
  285.5,     285.5,   285.5,   285.5,
  286.15,    286.15,  286.15,  286.15,
  286.6,     286.6,   286.6,   286.6,
  287.05,    287.05,  287.05,  287.05,
  287.7,     287.7,   287.7,   287.7,
  288.4,     288.4,   288.4,   288.4,
  288.95,    288.95,  288.95,  288.95,
  289.3,     289.3,   289.3,   289.3,
  289.3,     289.3,   289.3,   289.3,
  289,       289,     289,     289,
  289.05,    289.05,  289.05,  289.05,
  289.8,     289.8,   289.8,   289.8,
  290.45,    290.45,  290.45,  290.45,
  290.7,     290.7,   290.7,   290.7,
  290.85,    290.85,  290.85,  290.85,
  290.7,     290.7,   290.7,   290.7,
  290.3,     290.3,   290.3,   290.3,
  289.9,     289.9,   289.9,   289.9,
  289.95,    289.95,  289.95,  289.95,
  290.3,     290.3,   290.3,   290.3,
  290.5,     290.5,   290.5,   290.5,
  290.35,    290.35,  290.35,  290.35,
  290.2,     290.2,   290.2,   290.2,
  290.2,     290.2,   290.2,   290.2,
  290.1,     290.1,   290.1,   290.1,
  290.05,    290.05,  290.05,  290.05,
  290.1,     290.1,   290.1,   290.1,
  290.2,     290.2,   290.2,   290.2,
  290.15,    290.15,  290.15,  290.15,
  290.1,     290.1,   290.1,   290.1,
  290.25,    290.25,  290.25,  290.25,
  290.4,     290.4,   290.4,   290.4,
  290.4,     290.4,   290.4,   290.4,
  290.2,     290.2,   290.2,   290.2,
  290.1,     290.1,   290.1,   290.1,
  289.95,    289.95,  289.95,  289.95,
  289.55,    289.55,  289.55,  289.55,
  289.4,     289.4,   289.4,   289.4,
  289.4,     289.4,   289.4,   289.4,
  289.25,    289.25,  289.25,  289.25,
  289.15,    289.15,  289.15,  289.15,
  289.1,     289.1,   289.1,   289.1,
  289,       289,     289,     289,
  288.9,     288.9,   288.9,   288.9,
  288.8,     288.8,   288.8,   288.8,
  288.75,    288.75,  288.75,  288.75,
  288.8,     288.8,   288.8,   288.8,
  289,       289,     289,     289,
  289.45,    289.45,  289.45,  289.45,
  290.05,    290.05,  290.05,  290.05,
  290.55,    290.55,  290.55,  290.55,
  291,       291,     291,     291,
  291.5,     291.5,   291.5,   291.5,
  291.8,     291.8,   291.8,   291.8,
  292.05,    292.05,  292.05,  292.05,
  292.5,     292.5,   292.5,   292.5,
  292.75,    292.75,  292.75,  292.75,
  292.7,     292.7,   292.7,   292.7,
  292.95,    292.95,  292.95,  292.95,
  293.2,     293.2,   293.2,   293.2,
  293.45,    293.45,  293.45,  293.45,
  294.25,    294.25,  294.25,  294.25,
  294.95,    294.95,  294.95,  294.95,
  295.25,    295.25,  295.25,  295.25,
  295.15,    295.15,  295.15,  295.15,
  295,       295,     295,     295,
  295.2,     295.2,   295.2,   295.2,
  295.6,     295.6,   295.6,   295.6,
  295.8,     295.8,   295.8,   295.8,
  295.55,    295.55,  295.55,  295.55,
  295.05,    295.05,  295.05,  295.05,
  294.4,     294.4,   294.4,   294.4,
  293.65,    293.65,  293.65,  293.65,
  293.1,     293.1,   293.1,   293.1,
  293,       293,     293,     293,
  293.05,    293.05,  293.05,  293.05,
  292.95,    292.95,  292.95,  292.95,
  292.6,     292.6,   292.6,   292.6,
  292.3,     292.3,   292.3,   292.3,
  292.45,    292.45,  292.45,  292.45,
  292.7,     292.7,   292.7,   292.7,
  292.65,    292.65,  292.65,  292.65,
  292.45,    292.45,  292.45,  292.45,
  292.3,     292.3,   292.3,   292.3,
  292.2,     292.2,   292.2,   292.2,
  292.1,     292.1,   292.1,   292.1,
  291.9,     291.9,   291.9,   291.9,
  291.6,     291.6,   291.6,   291.6,
  291.25,    291.25,  291.25,  291.25,
  291,       291,     291,     291,
  290.85,    290.85,  290.85,  290.85,
  290.6,     290.6,   290.6,   290.6,
  290.4,     290.4,   290.4,   290.4,
  290.25,    290.25,  290.25,  290.25,
  290.15,    290.15,  290.15,  290.15,
  290.35,    290.35,  290.35,  290.35,
  290.95,    290.95,  290.95,  290.95,
  291.6,     291.6,   291.6,   291.6,
  292.05,    292.05,  292.05,  292.05,
  292.45,    292.45,  292.45,  292.45,
  292.95,    292.95,  292.95,  292.95,
  293.15,    293.15,  293.15,  293.15,
  293,       293,     293,     293,
  293.2,     293.2,   293.2,   293.2,
  293.55,    293.55,  293.55,  293.55,
  293.7,     293.7,   293.7,   293.7,
  294,       294,     294,     294,
  294.3,     294.3,   294.3,   294.3,
  294.3,     294.3,   294.3,   294.3,
  294.45,    294.45,  294.45,  294.45,
  294.8,     294.8,   294.8,   294.8,
  294.8,     294.8,   294.8,   294.8,
  294.55,    294.55,  294.55,  294.55,
  294.15,    294.15,  294.15,  294.15,
  293.75,    293.75,  293.75,  293.75,
  293.55,    293.55,  293.55,  293.55,
  293.25,    293.25,  293.25,  293.25,
  292.8,     292.8,   292.8,   292.8,
  292.3,     292.3,   292.3,   292.3,
  291.85,    291.85,  291.85,  291.85,
  291.25,    291.25,  291.25,  291.25,
  290.6,     290.6,   290.6,   290.6,
  290,       290,     290,     290,
  289.45,    289.45,  289.45,  289.45,
  289.15,    289.15,  289.15,  289.15,
  288.95,    288.95,  288.95,  288.95,
  288.8,     288.8,   288.8,   288.8,
  288.65,    288.65,  288.65,  288.65,
  288.45,    288.45,  288.45,  288.45,
  288.1,     288.1,   288.1,   288.1,
  287.6,     287.6,   287.6,   287.6,
  287.2,     287.2,   287.2,   287.2,
  287,       287,     287,     287,
  286.8,     286.8,   286.8,   286.8,
  286.35,    286.35,  286.35,  286.35,
  285.95,    285.95,  285.95,  285.95,
  285.7,     285.7,   285.7,   285.7,
  285.5,     285.5,   285.5,   285.5,
  285.5,     285.5,   285.5,   285.5,
  285.6,     285.6,   285.6,   285.6,
  285.7,     285.7,   285.7,   285.7,
  285.8,     285.8,   285.8,   285.8,
  285.9,     285.9,   285.9,   285.9,
  286.1,     286.1,   286.1,   286.1,
  286.35,    286.35,  286.35,  286.35,
  286.65,    286.65,  286.65,  286.65,
  286.95,    286.95,  286.95,  286.95,
  287.3,     287.3,   287.3,   287.3,
  287.7,     287.7,   287.7,   287.7,
  288,       288,     288,     288,
  288.4,     288.4,   288.4,   288.4,
  289,       289,     289,     289,
  289.85,    289.85,  289.85,  289.85,
  290.4,     290.4,   290.4,   290.4,
  290.8,     290.8,   290.8,   290.8,
  291.6,     291.6,   291.6,   291.6,
  292.4,     292.4,   292.4,   292.4,
  292.85,    292.85,  292.85,  292.85,
  293.15,    293.15,  293.15,  293.15,
  293.2,     293.2,   293.2,   293.2,
  293.3,     293.3,   293.3,   293.3,
  293.55,    293.55,  293.55,  293.55,
  293.4,     293.4,   293.4,   293.4,
  293.05,    293.05,  293.05,  293.05,
  292.55,    292.55,  292.55,  292.55,
  291.8,     291.8,   291.8,   291.8,
  291.2,     291.2,   291.2,   291.2,
  291,       291,     291,     291,
  290.6,     290.6,   290.6,   290.6,
  289.9,     289.9,   289.9,   289.9,
  289.35,    289.35,  289.35,  289.35,
  288.85,    288.85,  288.85,  288.85,
  288.4,     288.4,   288.4,   288.4,
  288.15,    288.15,  288.15,  288.15,
  287.95,    287.95,  287.95,  287.95,
  287.65,    287.65,  287.65,  287.65,
  287.35,    287.35,  287.35,  287.35,
  287.25,    287.25,  287.25,  287.25,
  286.9,     286.9,   286.9,   286.9,
  286.5,     286.5,   286.5,   286.5,
  286.25,    286.25,  286.25,  286.25,
  286.05,    286.05,  286.05,  286.05,
  285.8,     285.8,   285.8,   285.8,
  285.6,     285.6,   285.6,   285.6,
  285.6,     285.6,   285.6,   285.6,
  285.5,     285.5,   285.5,   285.5,
  285.35,    285.35,  285.35,  285.35,
  285.4,     285.4,   285.4,   285.4,
  285.35,    285.35,  285.35,  285.35,
  285.15,    285.15,  285.15,  285.15,
  285.05,    285.05,  285.05,  285.05,
  285.25,    285.25,  285.25,  285.25,
  285.9,     285.9,   285.9,   285.9,
  286.8,     286.8,   286.8,   286.8,
  288,       288,     288,     288,
  289.3,     289.3,   289.3,   289.3,
  290.5,     290.5,   290.5,   290.5,
  291.45,    291.45,  291.45,  291.45,
  292.25,    292.25,  292.25,  292.25,
  292.75,    292.75,  292.75,  292.75,
  293,       293,     293,     293,
  293.35,    293.35,  293.35,  293.35,
  293.6,     293.6,   293.6,   293.6,
  293.9,     293.9,   293.9,   293.9,
  294.3,     294.3,   294.3,   294.3,
  294.45,    294.45,  294.45,  294.45,
  294.25,    294.25,  294.25,  294.25,
  294.15,    294.15,  294.15,  294.15,
  294.25,    294.25,  294.25,  294.25,
  294.45,    294.45,  294.45,  294.45,
  294.45,    294.45,  294.45,  294.45,
  294.1,     294.1,   294.1,   294.1,
  293.8,     293.8,   293.8,   293.8,
  293.35,    293.35,  293.35,  293.35,
  293,       293,     293,     293,
  292.65,    292.65,  292.65,  292.65,
  291.85,    291.85,  291.85,  291.85,
  291,       291,     291,     291,
  290.45,    290.45,  290.45,  290.45,
  290.05,    290.05,  290.05,  290.05,
  289.8,     289.8,   289.8,   289.8,
  289.7,     289.7,   289.7,   289.7,
  289.55,    289.55,  289.55,  289.55,
  289.45,    289.45,  289.45,  289.45,
  289.4,     289.4,   289.4,   289.4,
  289.3,     289.3,   289.3,   289.3,
  289,       289,     289,     289,
  288.9,     288.9,   288.9,   288.9,
  288.8,     288.8,   288.8,   288.8,
  288.4,     288.4,   288.4,   288.4,
  288.25,    288.25,  288.25,  288.25,
  288.3,     288.3,   288.3,   288.3,
  288.3,     288.3,   288.3,   288.3,
  288.4,     288.4,   288.4,   288.4,
  288.6,     288.6,   288.6,   288.6,
  288.45,    288.45,  288.45,  288.45,
  288.25,    288.25,  288.25,  288.25,
  288.25,    288.25,  288.25,  288.25,
  288.25,    288.25,  288.25,  288.25,
  288.4,     288.4,   288.4,   288.4,
  288.65,    288.65,  288.65,  288.65,
  289.1,     289.1,   289.1,   289.1,
  289.9,     289.9,   289.9,   289.9,
  290.55,    290.55,  290.55,  290.55,
  290.85,    290.85,  290.85,  290.85,
  291,       291,     291,     291,
  291.6,     291.6,   291.6,   291.6,
  292.65,    292.65,  292.65,  292.65,
  293.65,    293.65,  293.65,  293.65,
  294.45,    294.45,  294.45,  294.45,
  294.8,     294.8,   294.8,   294.8,
  295.15,    295.15,  295.15,  295.15,
  295.65,    295.65,  295.65,  295.65,
  296.15,    296.15,  296.15,  296.15,
  296.35,    296.35,  296.35,  296.35,
  296.2,     296.2,   296.2,   296.2,
  296,       296,     296,     296,
  295.85,    295.85,  295.85,  295.85,
  295.75,    295.75,  295.75,  295.75,
  295.45,    295.45,  295.45,  295.45,
  295.15,    295.15,  295.15,  295.15,
  294.75,    294.75,  294.75,  294.75,
  294.1,     294.1,   294.1,   294.1,
  293.45,    293.45,  293.45,  293.45,
  292.85,    292.85,  292.85,  292.85,
  292.3,     292.3,   292.3,   292.3,
  291.95,    291.95,  291.95,  291.95,
  291.5,     291.5,   291.5,   291.5,
  291,       291,     291,     291,
  290.6,     290.6,   290.6,   290.6,
  289.85,    289.85,  289.85,  289.85,
  289.35,    289.35,  289.35,  289.35,
  289.45,    289.45,  289.45,  289.45,
  289.55,    289.55,  289.55,  289.55,
  289.5,     289.5,   289.5,   289.5,
  289.35,    289.35,  289.35,  289.35,
  289.3,     289.3,   289.3,   289.3,
  289.25,    289.25,  289.25,  289.25,
  289.05,    289.05,  289.05,  289.05,
  288.85,    288.85,  288.85,  288.85,
  288.75,    288.75,  288.75,  288.75,
  288.6,     288.6,   288.6,   288.6,
  288.25,    288.25,  288.25,  288.25,
  287.9,     287.9,   287.9,   287.9,
  287.65,    287.65,  287.65,  287.65,
  287.25,    287.25,  287.25,  287.25,
  286.85,    286.85,  286.85,  286.85,
  286.95,    286.95,  286.95,  286.95,
  287.45,    287.45,  287.45,  287.45,
  288.05,    288.05,  288.05,  288.05,
  288.45,    288.45,  288.45,  288.45,
  288.8,     288.8,   288.8,   288.8,
  289.55,    289.55,  289.55,  289.55,
  290.6,     290.6,   290.6,   290.6,
  291.25,    291.25,  291.25,  291.25,
  291.35,    291.35,  291.35,  291.35,
  291.35,    291.35,  291.35,  291.35,
  291.5,     291.5,   291.5,   291.5,
  291.7,     291.7,   291.7,   291.7,
  291.75,    291.75,  291.75,  291.75,
  291.95,    291.95,  291.95,  291.95,
  292.15,    292.15,  292.15,  292.15,
  292.3,     292.3,   292.3,   292.3,
  292.4,     292.4,   292.4,   292.4,
  292.35,    292.35,  292.35,  292.35,
  292.05,    292.05,  292.05,  292.05,
  291.8,     291.8,   291.8,   291.8,
  291.8,     291.8,   291.8,   291.8,
  291.55,    291.55,  291.55,  291.55,
  291.15,    291.15,  291.15,  291.15,
  290.75,    290.75,  290.75,  290.75,
  290.3,     290.3,   290.3,   290.3,
  289.95,    289.95,  289.95,  289.95,
  289.65,    289.65,  289.65,  289.65,
  289.35,    289.35,  289.35,  289.35,
  288.9,     288.9,   288.9,   288.9,
  288.2,     288.2,   288.2,   288.2,
  287.7,     287.7,   287.7,   287.7,
  287.5,     287.5,   287.5,   287.5,
  287.3,     287.3,   287.3,   287.3,
  286.7,     286.7,   286.7,   286.7,
  286.05,    286.05,  286.05,  286.05,
  285.8,     285.8,   285.8,   285.8,
  285.55,    285.55,  285.55,  285.55,
  285.25,    285.25,  285.25,  285.25,
  284.9,     284.9,   284.9,   284.9,
  284.5,     284.5,   284.5,   284.5,
  284.2,     284.2,   284.2,   284.2,
  284.1,     284.1,   284.1,   284.1,
  284.15,    284.15,  284.15,  284.15,
  284.05,    284.05,  284.05,  284.05,
  284.1,     284.1,   284.1,   284.1,
  284.15,    284.15,  284.15,  284.15,
  284.1,     284.1,   284.1,   284.1,
  284.3,     284.3,   284.3,   284.3,
  284.55,    284.55,  284.55,  284.55,
  285.35,    285.35,  285.35,  285.35,
  286.6,     286.6,   286.6,   286.6,
  287.7,     287.7,   287.7,   287.7,
  288.8,     288.8,   288.8,   288.8,
  289.65,    289.65,  289.65,  289.65,
  290.5,     290.5,   290.5,   290.5,
  290.9,     290.9,   290.9,   290.9,
  291,       291,     291,     291,
  291.2,     291.2,   291.2,   291.2,
  290.95,    290.95,  290.95,  290.95,
  291.3,     291.3,   291.3,   291.3,
  292.25,    292.25,  292.25,  292.25,
  292.6,     292.6,   292.6,   292.6,
  292.65,    292.65,  292.65,  292.65,
  292.65,    292.65,  292.65,  292.65,
  292.6,     292.6,   292.6,   292.6,
  292.5,     292.5,   292.5,   292.5,
  292.1,     292.1,   292.1,   292.1,
  291.7,     291.7,   291.7,   291.7,
  291.45,    291.45,  291.45,  291.45,
  291.2,     291.2,   291.2,   291.2,
  290.85,    290.85,  290.85,  290.85,
  290.15,    290.15,  290.15,  290.15,
  289.05,    289.05,  289.05,  289.05,
  288.2,     288.2,   288.2,   288.2,
  287.7,     287.7,   287.7,   287.7,
  287.15,    287.15,  287.15,  287.15,
  286.65,    286.65,  286.65,  286.65,
  286.3,     286.3,   286.3,   286.3,
  286.1,     286.1,   286.1,   286.1,
  286.2,     286.2,   286.2,   286.2,
  286.55,    286.55,  286.55,  286.55,
  287.1,     287.1,   287.1,   287.1,
  287.55,    287.55,  287.55,  287.55,
  287.2,     287.2,   287.2,   287.2,
  286.6,     286.6,   286.6,   286.6,
  286.4,     286.4,   286.4,   286.4,
  286.35,    286.35,  286.35,  286.35,
  286.35,    286.35,  286.35,  286.35,
  286.4,     286.4,   286.4,   286.4,
  286.4,     286.4,   286.4,   286.4,
  286.35,    286.35,  286.35,  286.35,
  286.35,    286.35,  286.35,  286.35,
  286.4,     286.4,   286.4,   286.4,
  286.45,    286.45,  286.45,  286.45,
  286.45,    286.45,  286.45,  286.45,
  286.45,    286.45,  286.45,  286.45,
  286.5,     286.5,   286.5,   286.5,
  286.65,    286.65,  286.65,  286.65,
  286.9,     286.9,   286.9,   286.9,
  287.1,     287.1,   287.1,   287.1,
  287.3,     287.3,   287.3,   287.3,
  287.65,    287.65,  287.65,  287.65,
  287.9,     287.9,   287.9,   287.9,
  288.2,     288.2,   288.2,   288.2,
  288.55,    288.55,  288.55,  288.55,
  288.2,     288.2,   288.2,   288.2,
  288.15,    288.15,  288.15,  288.15,
  288.95,    288.95,  288.95,  288.95,
  289.4,     289.4,   289.4,   289.4,
  290,       290,     290,     290,
  290.45,    290.45,  290.45,  290.45,
  290.5,     290.5,   290.5,   290.5,
  290.6,     290.6,   290.6,   290.6,
  290.8,     290.8,   290.8,   290.8,
  291.3,     291.3,   291.3,   291.3,
  291.35,    291.35,  291.35,  291.35,
  290.85,    290.85,  290.85,  290.85,
  290.5,     290.5,   290.5,   290.5,
  290.3,     290.3,   290.3,   290.3,
  289.8,     289.8,   289.8,   289.8,
  289.1,     289.1,   289.1,   289.1,
  288.45,    288.45,  288.45,  288.45,
  288.1,     288.1,   288.1,   288.1,
  287.95,    287.95,  287.95,  287.95,
  287.7,     287.7,   287.7,   287.7,
  287.1,     287.1,   287.1,   287.1,
  286.45,    286.45,  286.45,  286.45,
  286.15,    286.15,  286.15,  286.15,
  286,       286,     286,     286,
  286,       286,     286,     286,
  286,       286,     286,     286,
  286,       286,     286,     286,
  286.15,    286.15,  286.15,  286.15,
  286.3,     286.3,   286.3,   286.3,
  286.4,     286.4,   286.4,   286.4,
  286.55,    286.55,  286.55,  286.55,
  286.7,     286.7,   286.7,   286.7,
  286.8,     286.8,   286.8,   286.8,
  286.9,     286.9,   286.9,   286.9,
  287,       287,     287,     287,
  287.1,     287.1,   287.1,   287.1,
  287.2,     287.2,   287.2,   287.2,
  287.25,    287.25,  287.25,  287.25,
  287.3,     287.3,   287.3,   287.3,
  287.55,    287.55,  287.55,  287.55,
  288,       288,     288,     288,
  288.45,    288.45,  288.45,  288.45,
  288.9,     288.9,   288.9,   288.9,
  289.65,    289.65,  289.65,  289.65,
  290.35,    290.35,  290.35,  290.35,
  290.75,    290.75,  290.75,  290.75,
  290.9,     290.9,   290.9,   290.9,
  290.75,    290.75,  290.75,  290.75,
  290.45,    290.45,  290.45,  290.45,
  290.2,     290.2,   290.2,   290.2,
  290.2,     290.2,   290.2,   290.2,
  290.3,     290.3,   290.3,   290.3,
  290.45,    290.45,  290.45,  290.45,
  290.45,    290.45,  290.45,  290.45,
  290.35,    290.35,  290.35,  290.35,
  290.4,     290.4,   290.4,   290.4,
  290.35,    290.35,  290.35,  290.35,
  290.15,    290.15,  290.15,  290.15,
  289.9,     289.9,   289.9,   289.9,
  289.6,     289.6,   289.6,   289.6,
  289.3,     289.3,   289.3,   289.3,
  288.8,     288.8,   288.8,   288.8,
  288.4,     288.4,   288.4,   288.4,
  288.3,     288.3,   288.3,   288.3,
  288.25,    288.25,  288.25,  288.25,
  288.3,     288.3,   288.3,   288.3,
  288.35,    288.35,  288.35,  288.35,
  288.3,     288.3,   288.3,   288.3,
  288.2,     288.2,   288.2,   288.2,
  288.1,     288.1,   288.1,   288.1,
  288.05,    288.05,  288.05,  288.05,
  288.05,    288.05,  288.05,  288.05,
  287.9,     287.9,   287.9,   287.9,
  287.7,     287.7,   287.7,   287.7,
  287.65,    287.65,  287.65,  287.65,
  287.8,     287.8,   287.8,   287.8,
  287.75,    287.75,  287.75,  287.75,
  287.4,     287.4,   287.4,   287.4,
  287.1,     287.1,   287.1,   287.1,
  286.8,     286.8,   286.8,   286.8,
  286.6,     286.6,   286.6,   286.6,
  286.45,    286.45,  286.45,  286.45,
  286.25,    286.25,  286.25,  286.25,
  286.1,     286.1,   286.1,   286.1,
  286.15,    286.15,  286.15,  286.15,
  286.3,     286.3,   286.3,   286.3,
  286.55,    286.55,  286.55,  286.55,
  286.9,     286.9,   286.9,   286.9,
  287.3,     287.3,   287.3,   287.3,
  287.85,    287.85,  287.85,  287.85,
  288.4,     288.4,   288.4,   288.4,
  288.9,     288.9,   288.9,   288.9,
  289.25,    289.25,  289.25,  289.25,
  289.35,    289.35,  289.35,  289.35,
  289.65,    289.65,  289.65,  289.65,
  289.95,    289.95,  289.95,  289.95,
  290.2,     290.2,   290.2,   290.2,
  290.45,    290.45,  290.45,  290.45,
  290.6,     290.6,   290.6,   290.6,
  290.45,    290.45,  290.45,  290.45,
  290.25,    290.25,  290.25,  290.25,
  290.2,     290.2,   290.2,   290.2,
  290.05,    290.05,  290.05,  290.05,
  289.85,    289.85,  289.85,  289.85,
  289.35,    289.35,  289.35,  289.35,
  289.15,    289.15,  289.15,  289.15,
  289,       289,     289,     289,
  288.65,    288.65,  288.65,  288.65,
  288.5,     288.5,   288.5,   288.5,
  288.25,    288.25,  288.25,  288.25,
  287.75,    287.75,  287.75,  287.75,
  287.15,    287.15,  287.15,  287.15,
  286.8,     286.8,   286.8,   286.8,
  286.45,    286.45,  286.45,  286.45,
  285.85,    285.85,  285.85,  285.85,
  285.3,     285.3,   285.3,   285.3,
  284.8,     284.8,   284.8,   284.8,
  284.45,    284.45,  284.45,  284.45,
  284.4,     284.4,   284.4,   284.4,
  284.55,    284.55,  284.55,  284.55,
  284.95,    284.95,  284.95,  284.95,
  285.3,     285.3,   285.3,   285.3,
  285.35,    285.35,  285.35,  285.35,
  285.25,    285.25,  285.25,  285.25,
  285.1,     285.1,   285.1,   285.1,
  284.95,    284.95,  284.95,  284.95,
  284.6,     284.6,   284.6,   284.6,
  284.15,    284.15,  284.15,  284.15,
  283.75,    283.75,  283.75,  283.75,
  283.45,    283.45,  283.45,  283.45,
  283.3,     283.3,   283.3,   283.3,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.35,    283.35,  283.35,  283.35,
  283.5,     283.5,   283.5,   283.5,
  283.65,    283.65,  283.65,  283.65,
  283.95,    283.95,  283.95,  283.95,
  284.9,     284.9,   284.9,   284.9,
  285.75,    285.75,  285.75,  285.75,
  286.35,    286.35,  286.35,  286.35,
  287.2,     287.2,   287.2,   287.2,
  287.5,     287.5,   287.5,   287.5,
  287.6,     287.6,   287.6,   287.6,
  287.85,    287.85,  287.85,  287.85,
  288.05,    288.05,  288.05,  288.05,
  288.2,     288.2,   288.2,   288.2,
  288.3,     288.3,   288.3,   288.3,
  288.45,    288.45,  288.45,  288.45,
  288.7,     288.7,   288.7,   288.7,
  289.15,    289.15,  289.15,  289.15,
  289.3,     289.3,   289.3,   289.3,
  289.35,    289.35,  289.35,  289.35,
  289.6,     289.6,   289.6,   289.6,
  289.6,     289.6,   289.6,   289.6,
  289.15,    289.15,  289.15,  289.15,
  288.8,     288.8,   288.8,   288.8,
  288.75,    288.75,  288.75,  288.75,
  288.4,     288.4,   288.4,   288.4,
  287.7,     287.7,   287.7,   287.7,
  287.1,     287.1,   287.1,   287.1,
  286.6,     286.6,   286.6,   286.6,
  285.95,    285.95,  285.95,  285.95,
  285.35,    285.35,  285.35,  285.35,
  284.95,    284.95,  284.95,  284.95,
  284.65,    284.65,  284.65,  284.65,
  284.2,     284.2,   284.2,   284.2,
  283.95,    283.95,  283.95,  283.95,
  283.75,    283.75,  283.75,  283.75,
  283.15,    283.15,  283.15,  283.15,
  282.1,     282.1,   282.1,   282.1,
  281.55,    281.55,  281.55,  281.55,
  281.65,    281.65,  281.65,  281.65,
  281.45,    281.45,  281.45,  281.45,
  281.35,    281.35,  281.35,  281.35,
  281.5,     281.5,   281.5,   281.5,
  281.5,     281.5,   281.5,   281.5,
  281.65,    281.65,  281.65,  281.65,
  281.65,    281.65,  281.65,  281.65,
  281.25,    281.25,  281.25,  281.25,
  281.05,    281.05,  281.05,  281.05,
  281,       281,     281,     281,
  281.15,    281.15,  281.15,  281.15,
  281.4,     281.4,   281.4,   281.4,
  281.85,    281.85,  281.85,  281.85,
  282.75,    282.75,  282.75,  282.75,
  283.75,    283.75,  283.75,  283.75,
  284.9,     284.9,   284.9,   284.9,
  286.3,     286.3,   286.3,   286.3,
  287.65,    287.65,  287.65,  287.65,
  288.45,    288.45,  288.45,  288.45,
  288.9,     288.9,   288.9,   288.9,
  289.45,    289.45,  289.45,  289.45,
  289.95,    289.95,  289.95,  289.95,
  290.25,    290.25,  290.25,  290.25,
  290.5,     290.5,   290.5,   290.5,
  290.85,    290.85,  290.85,  290.85,
  291.2,     291.2,   291.2,   291.2,
  291.5,     291.5,   291.5,   291.5,
  291.5,     291.5,   291.5,   291.5,
  291.3,     291.3,   291.3,   291.3,
  291.25,    291.25,  291.25,  291.25,
  291.15,    291.15,  291.15,  291.15,
  291,       291,     291,     291,
  290.8,     290.8,   290.8,   290.8,
  290.7,     290.7,   290.7,   290.7,
  290.65,    290.65,  290.65,  290.65,
  290.3,     290.3,   290.3,   290.3,
  289.6,     289.6,   289.6,   289.6,
  288.8,     288.8,   288.8,   288.8,
  288.2,     288.2,   288.2,   288.2,
  287.6,     287.6,   287.6,   287.6,
  287.1,     287.1,   287.1,   287.1,
  287.05,    287.05,  287.05,  287.05,
  287.3,     287.3,   287.3,   287.3,
  287.4,     287.4,   287.4,   287.4,
  287.35,    287.35,  287.35,  287.35,
  287.6,     287.6,   287.6,   287.6,
  287.8,     287.8,   287.8,   287.8,
  287.9,     287.9,   287.9,   287.9,
  288.05,    288.05,  288.05,  288.05,
  288,       288,     288,     288,
  288.05,    288.05,  288.05,  288.05,
  288.2,     288.2,   288.2,   288.2,
  288.15,    288.15,  288.15,  288.15,
  287.95,    287.95,  287.95,  287.95,
  287.55,    287.55,  287.55,  287.55,
  287.2,     287.2,   287.2,   287.2,
  287.25,    287.25,  287.25,  287.25,
  287.5,     287.5,   287.5,   287.5,
  287.75,    287.75,  287.75,  287.75,
  287.9,     287.9,   287.9,   287.9,
  288,       288,     288,     288,
  288.25,    288.25,  288.25,  288.25,
  288.7,     288.7,   288.7,   288.7,
  289.1,     289.1,   289.1,   289.1,
  289.35,    289.35,  289.35,  289.35,
  289.5,     289.5,   289.5,   289.5,
  289.7,     289.7,   289.7,   289.7,
  290.15,    290.15,  290.15,  290.15,
  290.5,     290.5,   290.5,   290.5,
  290.8,     290.8,   290.8,   290.8,
  291.15,    291.15,  291.15,  291.15,
  291.05,    291.05,  291.05,  291.05,
  291,       291,     291,     291,
  291.45,    291.45,  291.45,  291.45,
  291.6,     291.6,   291.6,   291.6,
  291.4,     291.4,   291.4,   291.4,
  291.25,    291.25,  291.25,  291.25,
  291.05,    291.05,  291.05,  291.05,
  290.9,     290.9,   290.9,   290.9,
  290.9,     290.9,   290.9,   290.9,
  290.95,    290.95,  290.95,  290.95,
  290.95,    290.95,  290.95,  290.95,
  290.95,    290.95,  290.95,  290.95,
  290.85,    290.85,  290.85,  290.85,
  290.65,    290.65,  290.65,  290.65,
  290.45,    290.45,  290.45,  290.45,
  288.85,    288.85,  288.85,  288.85,
  287.2,     287.2,   287.2,   287.2,
  286.9,     286.9,   286.9,   286.9,
  286.5,     286.5,   286.5,   286.5,
  286.15,    286.15,  286.15,  286.15,
  286,       286,     286,     286,
  285.85,    285.85,  285.85,  285.85,
  285.65,    285.65,  285.65,  285.65,
  285.45,    285.45,  285.45,  285.45,
  285.15,    285.15,  285.15,  285.15,
  284.9,     284.9,   284.9,   284.9,
  285,       285,     285,     285,
  285.3,     285.3,   285.3,   285.3,
  285.25,    285.25,  285.25,  285.25,
  284.9,     284.9,   284.9,   284.9,
  284.7,     284.7,   284.7,   284.7,
  284.4,     284.4,   284.4,   284.4,
  283.9,     283.9,   283.9,   283.9,
  283.4,     283.4,   283.4,   283.4,
  282.9,     282.9,   282.9,   282.9,
  282.55,    282.55,  282.55,  282.55,
  282.5,     282.5,   282.5,   282.5,
  282.8,     282.8,   282.8,   282.8,
  283.5,     283.5,   283.5,   283.5,
  284.3,     284.3,   284.3,   284.3,
  284.7,     284.7,   284.7,   284.7,
  285.4,     285.4,   285.4,   285.4,
  286.35,    286.35,  286.35,  286.35,
  286.45,    286.45,  286.45,  286.45,
  286.95,    286.95,  286.95,  286.95,
  287.8,     287.8,   287.8,   287.8,
  287.95,    287.95,  287.95,  287.95,
  287.9,     287.9,   287.9,   287.9,
  287.8,     287.8,   287.8,   287.8,
  287.85,    287.85,  287.85,  287.85,
  288.05,    288.05,  288.05,  288.05,
  288.1,     288.1,   288.1,   288.1,
  288.05,    288.05,  288.05,  288.05,
  288,       288,     288,     288,
  288.05,    288.05,  288.05,  288.05,
  286.9,     286.9,   286.9,   286.9,
  285.05,    285.05,  285.05,  285.05,
  284.8,     284.8,   284.8,   284.8,
  285.3,     285.3,   285.3,   285.3,
  285.35,    285.35,  285.35,  285.35,
  284.75,    284.75,  284.75,  284.75,
  283.7,     283.7,   283.7,   283.7,
  282.85,    282.85,  282.85,  282.85,
  282.5,     282.5,   282.5,   282.5,
  282.7,     282.7,   282.7,   282.7,
  282.7,     282.7,   282.7,   282.7,
  282.05,    282.05,  282.05,  282.05,
  282.1,     282.1,   282.1,   282.1,
  282.95,    282.95,  282.95,  282.95,
  282.95,    282.95,  282.95,  282.95,
  282.3,     282.3,   282.3,   282.3,
  282.05,    282.05,  282.05,  282.05,
  282.1,     282.1,   282.1,   282.1,
  282.15,    282.15,  282.15,  282.15,
  282.2,     282.2,   282.2,   282.2,
  282.45,    282.45,  282.45,  282.45,
  282.45,    282.45,  282.45,  282.45,
  282.2,     282.2,   282.2,   282.2,
  282.15,    282.15,  282.15,  282.15,
  282.15,    282.15,  282.15,  282.15,
  282.25,    282.25,  282.25,  282.25,
  282.15,    282.15,  282.15,  282.15,
  281.6,     281.6,   281.6,   281.6,
  280.95,    280.95,  280.95,  280.95,
  280.9,     280.9,   280.9,   280.9,
  281.2,     281.2,   281.2,   281.2,
  281.85,    281.85,  281.85,  281.85,
  283.25,    283.25,  283.25,  283.25,
  284.7,     284.7,   284.7,   284.7,
  285.8,     285.8,   285.8,   285.8,
  286.75,    286.75,  286.75,  286.75,
  287.5,     287.5,   287.5,   287.5,
  287.6,     287.6,   287.6,   287.6,
  288,       288,     288,     288,
  288.75,    288.75,  288.75,  288.75,
  289.05,    289.05,  289.05,  289.05,
  288.85,    288.85,  288.85,  288.85,
  288.7,     288.7,   288.7,   288.7,
  288.8,     288.8,   288.8,   288.8,
  288.75,    288.75,  288.75,  288.75,
  288.7,     288.7,   288.7,   288.7,
  288.65,    288.65,  288.65,  288.65,
  288.9,     288.9,   288.9,   288.9,
  289.2,     289.2,   289.2,   289.2,
  289,       289,     289,     289,
  288.65,    288.65,  288.65,  288.65,
  288.3,     288.3,   288.3,   288.3,
  287.95,    287.95,  287.95,  287.95,
  287.4,     287.4,   287.4,   287.4,
  286.45,    286.45,  286.45,  286.45,
  285.55,    285.55,  285.55,  285.55,
  284.9,     284.9,   284.9,   284.9,
  284.5,     284.5,   284.5,   284.5,
  284.15,    284.15,  284.15,  284.15,
  283.7,     283.7,   283.7,   283.7,
  283.4,     283.4,   283.4,   283.4,
  283.3,     283.3,   283.3,   283.3,
  283.1,     283.1,   283.1,   283.1,
  282.7,     282.7,   282.7,   282.7,
  282.4,     282.4,   282.4,   282.4,
  282.25,    282.25,  282.25,  282.25,
  282.2,     282.2,   282.2,   282.2,
  282.3,     282.3,   282.3,   282.3,
  282.3,     282.3,   282.3,   282.3,
  282.15,    282.15,  282.15,  282.15,
  281.55,    281.55,  281.55,  281.55,
  280.9,     280.9,   280.9,   280.9,
  280.85,    280.85,  280.85,  280.85,
  281.05,    281.05,  281.05,  281.05,
  281.2,     281.2,   281.2,   281.2,
  281.4,     281.4,   281.4,   281.4,
  281.8,     281.8,   281.8,   281.8,
  282.1,     282.1,   282.1,   282.1,
  282.4,     282.4,   282.4,   282.4,
  283.1,     283.1,   283.1,   283.1,
  284,       284,     284,     284,
  285,       285,     285,     285,
  286.05,    286.05,  286.05,  286.05,
  287.05,    287.05,  287.05,  287.05,
  287.8,     287.8,   287.8,   287.8,
  288.2,     288.2,   288.2,   288.2,
  288.45,    288.45,  288.45,  288.45,
  288.9,     288.9,   288.9,   288.9,
  289.4,     289.4,   289.4,   289.4,
  289.6,     289.6,   289.6,   289.6,
  289.75,    289.75,  289.75,  289.75,
  289.95,    289.95,  289.95,  289.95,
  290.2,     290.2,   290.2,   290.2,
  290.45,    290.45,  290.45,  290.45,
  290.45,    290.45,  290.45,  290.45,
  290.4,     290.4,   290.4,   290.4,
  290.55,    290.55,  290.55,  290.55,
  290.55,    290.55,  290.55,  290.55,
  290.3,     290.3,   290.3,   290.3,
  290,       290,     290,     290,
  289.6,     289.6,   289.6,   289.6,
  288.9,     288.9,   288.9,   288.9,
  287.95,    287.95,  287.95,  287.95,
  287.1,     287.1,   287.1,   287.1,
  286.5,     286.5,   286.5,   286.5,
  285.95,    285.95,  285.95,  285.95,
  285.6,     285.6,   285.6,   285.6,
  285.35,    285.35,  285.35,  285.35,
  285,       285,     285,     285,
  284.9,     284.9,   284.9,   284.9,
  284.75,    284.75,  284.75,  284.75,
  284.65,    284.65,  284.65,  284.65,
  284.75,    284.75,  284.75,  284.75,
  284.95,    284.95,  284.95,  284.95,
  285,       285,     285,     285,
  284.65,    284.65,  284.65,  284.65,
  284.4,     284.4,   284.4,   284.4,
  284,       284,     284,     284,
  283.5,     283.5,   283.5,   283.5,
  283.5,     283.5,   283.5,   283.5,
  283.75,    283.75,  283.75,  283.75,
  283.35,    283.35,  283.35,  283.35,
  282.55,    282.55,  282.55,  282.55,
  282,       282,     282,     282,
  281.55,    281.55,  281.55,  281.55,
  281.4,     281.4,   281.4,   281.4,
  281.8,     281.8,   281.8,   281.8,
  282.85,    282.85,  282.85,  282.85,
  284.3,     284.3,   284.3,   284.3,
  286,       286,     286,     286,
  287.55,    287.55,  287.55,  287.55,
  288.55,    288.55,  288.55,  288.55,
  289.35,    289.35,  289.35,  289.35,
  289.95,    289.95,  289.95,  289.95,
  290.7,     290.7,   290.7,   290.7,
  291.35,    291.35,  291.35,  291.35,
  291.8,     291.8,   291.8,   291.8,
  292.4,     292.4,   292.4,   292.4,
  292.9,     292.9,   292.9,   292.9,
  293.3,     293.3,   293.3,   293.3,
  293.7,     293.7,   293.7,   293.7,
  294,       294,     294,     294,
  294.25,    294.25,  294.25,  294.25,
  294.55,    294.55,  294.55,  294.55,
  294.6,     294.6,   294.6,   294.6,
  294.35,    294.35,  294.35,  294.35,
  293.85,    293.85,  293.85,  293.85,
  293.05,    293.05,  293.05,  293.05,
  292.1,     292.1,   292.1,   292.1,
  291.25,    291.25,  291.25,  291.25,
  290.4,     290.4,   290.4,   290.4,
  289.7,     289.7,   289.7,   289.7,
  289.2,     289.2,   289.2,   289.2,
  288.75,    288.75,  288.75,  288.75,
  288.4,     288.4,   288.4,   288.4,
  288.15,    288.15,  288.15,  288.15,
  287.95,    287.95,  287.95,  287.95,
  287.9,     287.9,   287.9,   287.9,
  288.1,     288.1,   288.1,   288.1,
  288.45,    288.45,  288.45,  288.45,
  288.5,     288.5,   288.5,   288.5,
  287.95,    287.95,  287.95,  287.95,
  287.15,    287.15,  287.15,  287.15,
  286.6,     286.6,   286.6,   286.6,
  286.2,     286.2,   286.2,   286.2,
  285.85,    285.85,  285.85,  285.85,
  285.8,     285.8,   285.8,   285.8,
  285.65,    285.65,  285.65,  285.65,
  285.35,    285.35,  285.35,  285.35,
  285.1,     285.1,   285.1,   285.1,
  284.9,     284.9,   284.9,   284.9,
  284.8,     284.8,   284.8,   284.8,
  284.75,    284.75,  284.75,  284.75,
  284.75,    284.75,  284.75,  284.75,
  284.7,     284.7,   284.7,   284.7,
  284.9,     284.9,   284.9,   284.9,
  285.75,    285.75,  285.75,  285.75,
  286.85,    286.85,  286.85,  286.85,
  287.9,     287.9,   287.9,   287.9,
  288.85,    288.85,  288.85,  288.85,
  289.7,     289.7,   289.7,   289.7,
  290.4,     290.4,   290.4,   290.4,
  290.8,     290.8,   290.8,   290.8,
  290.8,     290.8,   290.8,   290.8,
  290.7,     290.7,   290.7,   290.7,
  290.7,     290.7,   290.7,   290.7,
  290.75,    290.75,  290.75,  290.75,
  290.85,    290.85,  290.85,  290.85,
  290.9,     290.9,   290.9,   290.9,
  291,       291,     291,     291,
  291,       291,     291,     291,
  290.7,     290.7,   290.7,   290.7,
  290.55,    290.55,  290.55,  290.55,
  290.4,     290.4,   290.4,   290.4,
  290.05,    290.05,  290.05,  290.05,
  289.95,    289.95,  289.95,  289.95,
  289.9,     289.9,   289.9,   289.9,
  289.75,    289.75,  289.75,  289.75,
  289.55,    289.55,  289.55,  289.55,
  289.35,    289.35,  289.35,  289.35,
  289.2,     289.2,   289.2,   289.2,
  289.1,     289.1,   289.1,   289.1,
  288.95,    288.95,  288.95,  288.95,
  288.7,     288.7,   288.7,   288.7,
  288.35,    288.35,  288.35,  288.35,
  287.9,     287.9,   287.9,   287.9,
  287.4,     287.4,   287.4,   287.4,
  286.95,    286.95,  286.95,  286.95,
  286.45,    286.45,  286.45,  286.45,
  286,       286,     286,     286,
  285.7,     285.7,   285.7,   285.7,
  285.4,     285.4,   285.4,   285.4,
  285.25,    285.25,  285.25,  285.25,
  285.15,    285.15,  285.15,  285.15,
  284.95,    284.95,  284.95,  284.95,
  284.75,    284.75,  284.75,  284.75,
  284.55,    284.55,  284.55,  284.55,
  284.45,    284.45,  284.45,  284.45,
  284.45,    284.45,  284.45,  284.45,
  284.45,    284.45,  284.45,  284.45,
  284.45,    284.45,  284.45,  284.45,
  284.6,     284.6,   284.6,   284.6,
  284.85,    284.85,  284.85,  284.85,
  285.3,     285.3,   285.3,   285.3,
  285.95,    285.95,  285.95,  285.95,
  286.65,    286.65,  286.65,  286.65,
  287.4,     287.4,   287.4,   287.4,
  288.3,     288.3,   288.3,   288.3,
  289.35,    289.35,  289.35,  289.35,
  290.15,    290.15,  290.15,  290.15,
  290.85,    290.85,  290.85,  290.85,
  291.3,     291.3,   291.3,   291.3,
  291.7,     291.7,   291.7,   291.7,
  292.4,     292.4,   292.4,   292.4,
  292.95,    292.95,  292.95,  292.95,
  293.25,    293.25,  293.25,  293.25,
  293.45,    293.45,  293.45,  293.45,
  293.5,     293.5,   293.5,   293.5,
  293.5,     293.5,   293.5,   293.5,
  293.4,     293.4,   293.4,   293.4,
  293.1,     293.1,   293.1,   293.1,
  292.8,     292.8,   292.8,   292.8,
  292.35,    292.35,  292.35,  292.35,
  291.8,     291.8,   291.8,   291.8,
  291.25,    291.25,  291.25,  291.25,
  290.4,     290.4,   290.4,   290.4,
  289.4,     289.4,   289.4,   289.4,
  288.5,     288.5,   288.5,   288.5,
  287.75,    287.75,  287.75,  287.75,
  287.2,     287.2,   287.2,   287.2,
  286.6,     286.6,   286.6,   286.6,
  286.15,    286.15,  286.15,  286.15,
  285.9,     285.9,   285.9,   285.9,
  285.55,    285.55,  285.55,  285.55,
  285.35,    285.35,  285.35,  285.35,
  285.25,    285.25,  285.25,  285.25,
  285.4,     285.4,   285.4,   285.4,
  285.8,     285.8,   285.8,   285.8,
  285.95,    285.95,  285.95,  285.95,
  285.9,     285.9,   285.9,   285.9,
  285.85,    285.85,  285.85,  285.85,
  285.7,     285.7,   285.7,   285.7,
  285.45,    285.45,  285.45,  285.45,
  285.3,     285.3,   285.3,   285.3,
  285.2,     285.2,   285.2,   285.2,
  285,       285,     285,     285,
  284.7,     284.7,   284.7,   284.7,
  284.45,    284.45,  284.45,  284.45,
  284.3,     284.3,   284.3,   284.3,
  284.35,    284.35,  284.35,  284.35,
  284.6,     284.6,   284.6,   284.6,
  284.9,     284.9,   284.9,   284.9,
  285.2,     285.2,   285.2,   285.2,
  285.55,    285.55,  285.55,  285.55,
  286.1,     286.1,   286.1,   286.1,
  286.85,    286.85,  286.85,  286.85,
  287.7,     287.7,   287.7,   287.7,
  288.35,    288.35,  288.35,  288.35,
  288.6,     288.6,   288.6,   288.6,
  289.05,    289.05,  289.05,  289.05,
  289.55,    289.55,  289.55,  289.55,
  289.6,     289.6,   289.6,   289.6,
  289.7,     289.7,   289.7,   289.7,
  289.65,    289.65,  289.65,  289.65,
  289.3,     289.3,   289.3,   289.3,
  289.4,     289.4,   289.4,   289.4,
  289.8,     289.8,   289.8,   289.8,
  289.9,     289.9,   289.9,   289.9,
  289.7,     289.7,   289.7,   289.7,
  289.3,     289.3,   289.3,   289.3,
  288.8,     288.8,   288.8,   288.8,
  288.25,    288.25,  288.25,  288.25,
  287.55,    287.55,  287.55,  287.55,
  286.75,    286.75,  286.75,  286.75,
  285.85,    285.85,  285.85,  285.85,
  284.75,    284.75,  284.75,  284.75,
  283.85,    283.85,  283.85,  283.85,
  283.4,     283.4,   283.4,   283.4,
  283,       283,     283,     283,
  282.7,     282.7,   282.7,   282.7,
  282.45,    282.45,  282.45,  282.45,
  282.1,     282.1,   282.1,   282.1,
  281.95,    281.95,  281.95,  281.95,
  281.75,    281.75,  281.75,  281.75,
  281.4,     281.4,   281.4,   281.4,
  281,       281,     281,     281,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.45,    280.45,  280.45,  280.45,
  280.1,     280.1,   280.1,   280.1,
  279.8,     279.8,   279.8,   279.8,
  279.6,     279.6,   279.6,   279.6,
  279.5,     279.5,   279.5,   279.5,
  279.05,    279.05,  279.05,  279.05,
  278.3,     278.3,   278.3,   278.3,
  277.7,     277.7,   277.7,   277.7,
  277.6,     277.6,   277.6,   277.6,
  277.65,    277.65,  277.65,  277.65,
  277.6,     277.6,   277.6,   277.6,
  278.5,     278.5,   278.5,   278.5,
  280.4,     280.4,   280.4,   280.4,
  282.35,    282.35,  282.35,  282.35,
  284.1,     284.1,   284.1,   284.1,
  285.5,     285.5,   285.5,   285.5,
  286.15,    286.15,  286.15,  286.15,
  286.4,     286.4,   286.4,   286.4,
  286.6,     286.6,   286.6,   286.6,
  286.85,    286.85,  286.85,  286.85,
  287.15,    287.15,  287.15,  287.15,
  287.2,     287.2,   287.2,   287.2,
  287.05,    287.05,  287.05,  287.05,
  287.45,    287.45,  287.45,  287.45,
  287.85,    287.85,  287.85,  287.85,
  287.9,     287.9,   287.9,   287.9,
  287.95,    287.95,  287.95,  287.95,
  288.05,    288.05,  288.05,  288.05,
  288.2,     288.2,   288.2,   288.2,
  288.1,     288.1,   288.1,   288.1,
  288,       288,     288,     288,
  287.3,     287.3,   287.3,   287.3,
  286.3,     286.3,   286.3,   286.3,
  285.65,    285.65,  285.65,  285.65,
  284.95,    284.95,  284.95,  284.95,
  284.15,    284.15,  284.15,  284.15,
  283.4,     283.4,   283.4,   283.4,
  282.8,     282.8,   282.8,   282.8,
  282.65,    282.65,  282.65,  282.65,
  282.75,    282.75,  282.75,  282.75,
  282.5,     282.5,   282.5,   282.5,
  282.15,    282.15,  282.15,  282.15,
  282,       282,     282,     282,
  281.8,     281.8,   281.8,   281.8,
  281.55,    281.55,  281.55,  281.55,
  281.35,    281.35,  281.35,  281.35,
  281.05,    281.05,  281.05,  281.05,
  280.65,    280.65,  280.65,  280.65,
  280.4,     280.4,   280.4,   280.4,
  280.2,     280.2,   280.2,   280.2,
  279.9,     279.9,   279.9,   279.9,
  279.7,     279.7,   279.7,   279.7,
  279.6,     279.6,   279.6,   279.6,
  279.55,    279.55,  279.55,  279.55,
  279.5,     279.5,   279.5,   279.5,
  279.4,     279.4,   279.4,   279.4,
  279.25,    279.25,  279.25,  279.25,
  279.2,     279.2,   279.2,   279.2,
  279.6,     279.6,   279.6,   279.6,
  280.5,     280.5,   280.5,   280.5,
  281.7,     281.7,   281.7,   281.7,
  282.8,     282.8,   282.8,   282.8,
  283.7,     283.7,   283.7,   283.7,
  284.5,     284.5,   284.5,   284.5,
  285.4,     285.4,   285.4,   285.4,
  286.25,    286.25,  286.25,  286.25,
  286.7,     286.7,   286.7,   286.7,
  286.95,    286.95,  286.95,  286.95,
  287.35,    287.35,  287.35,  287.35,
  287.7,     287.7,   287.7,   287.7,
  287.95,    287.95,  287.95,  287.95,
  288.25,    288.25,  288.25,  288.25,
  288.4,     288.4,   288.4,   288.4,
  288.55,    288.55,  288.55,  288.55,
  288.75,    288.75,  288.75,  288.75,
  288.8,     288.8,   288.8,   288.8,
  288.85,    288.85,  288.85,  288.85,
  288.85,    288.85,  288.85,  288.85,
  288.65,    288.65,  288.65,  288.65,
  288.35,    288.35,  288.35,  288.35,
  287.8,     287.8,   287.8,   287.8,
  287,       287,     287,     287,
  286.05,    286.05,  286.05,  286.05,
  285.1,     285.1,   285.1,   285.1,
  284.35,    284.35,  284.35,  284.35,
  283.75,    283.75,  283.75,  283.75,
  283.2,     283.2,   283.2,   283.2,
  282.75,    282.75,  282.75,  282.75,
  282.5,     282.5,   282.5,   282.5,
  282.35,    282.35,  282.35,  282.35,
  282.25,    282.25,  282.25,  282.25,
  282.15,    282.15,  282.15,  282.15,
  281.85,    281.85,  281.85,  281.85,
  281.4,     281.4,   281.4,   281.4,
  281.1,     281.1,   281.1,   281.1,
  281.05,    281.05,  281.05,  281.05,
  281.05,    281.05,  281.05,  281.05,
  281,       281,     281,     281,
  280.95,    280.95,  280.95,  280.95,
  280.85,    280.85,  280.85,  280.85,
  280.6,     280.6,   280.6,   280.6,
  280.35,    280.35,  280.35,  280.35,
  280.1,     280.1,   280.1,   280.1,
  279.8,     279.8,   279.8,   279.8,
  279.55,    279.55,  279.55,  279.55,
  279.4,     279.4,   279.4,   279.4,
  279.75,    279.75,  279.75,  279.75,
  280.75,    280.75,  280.75,  280.75,
  281.85,    281.85,  281.85,  281.85,
  283,       283,     283,     283,
  284.3,     284.3,   284.3,   284.3,
  285.6,     285.6,   285.6,   285.6,
  286.9,     286.9,   286.9,   286.9,
  287.9,     287.9,   287.9,   287.9,
  288.5,     288.5,   288.5,   288.5,
  288.95,    288.95,  288.95,  288.95,
  289.35,    289.35,  289.35,  289.35,
  289.8,     289.8,   289.8,   289.8,
  290.25,    290.25,  290.25,  290.25,
  290.65,    290.65,  290.65,  290.65,
  291.15,    291.15,  291.15,  291.15,
  291.5,     291.5,   291.5,   291.5,
  291.55,    291.55,  291.55,  291.55,
  291.55,    291.55,  291.55,  291.55,
  291.45,    291.45,  291.45,  291.45,
  291.25,    291.25,  291.25,  291.25,
  290.95,    290.95,  290.95,  290.95,
  290.5,     290.5,   290.5,   290.5,
  289.75,    289.75,  289.75,  289.75,
  288.75,    288.75,  288.75,  288.75,
  287.75,    287.75,  287.75,  287.75,
  286.7,     286.7,   286.7,   286.7,
  285.8,     285.8,   285.8,   285.8,
  285.25,    285.25,  285.25,  285.25,
  284.75,    284.75,  284.75,  284.75,
  284.1,     284.1,   284.1,   284.1,
  283.7,     283.7,   283.7,   283.7,
  283.6,     283.6,   283.6,   283.6,
  283.2,     283.2,   283.2,   283.2,
  282.7,     282.7,   282.7,   282.7,
  282.5,     282.5,   282.5,   282.5,
  282.6,     282.6,   282.6,   282.6,
  282.85,    282.85,  282.85,  282.85,
  282.95,    282.95,  282.95,  282.95,
  282.85,    282.85,  282.85,  282.85,
  282.65,    282.65,  282.65,  282.65,
  282.4,     282.4,   282.4,   282.4,
  282,       282,     282,     282,
  281.45,    281.45,  281.45,  281.45,
  281.1,     281.1,   281.1,   281.1,
  281,       281,     281,     281,
  280.95,    280.95,  280.95,  280.95,
  280.8,     280.8,   280.8,   280.8,
  280.65,    280.65,  280.65,  280.65,
  280.95,    280.95,  280.95,  280.95,
  281.5,     281.5,   281.5,   281.5,
  282.4,     282.4,   282.4,   282.4,
  283.95,    283.95,  283.95,  283.95,
  285.55,    285.55,  285.55,  285.55,
  286.9,     286.9,   286.9,   286.9,
  287.7,     287.7,   287.7,   287.7,
  287.9,     287.9,   287.9,   287.9,
  288.2,     288.2,   288.2,   288.2,
  288.6,     288.6,   288.6,   288.6,
  288.8,     288.8,   288.8,   288.8,
  289.05,    289.05,  289.05,  289.05,
  289.45,    289.45,  289.45,  289.45,
  289.75,    289.75,  289.75,  289.75,
  289.95,    289.95,  289.95,  289.95,
  290.05,    290.05,  290.05,  290.05,
  289.85,    289.85,  289.85,  289.85,
  289.35,    289.35,  289.35,  289.35,
  288.75,    288.75,  288.75,  288.75,
  288.25,    288.25,  288.25,  288.25,
  287.95,    287.95,  287.95,  287.95,
  287.75,    287.75,  287.75,  287.75,
  287.55,    287.55,  287.55,  287.55,
  287.3,     287.3,   287.3,   287.3,
  286.95,    286.95,  286.95,  286.95,
  286.5,     286.5,   286.5,   286.5,
  286.2,     286.2,   286.2,   286.2,
  286.1,     286.1,   286.1,   286.1,
  286,       286,     286,     286,
  286,       286,     286,     286,
  286.05,    286.05,  286.05,  286.05,
  286,       286,     286,     286,
  285.85,    285.85,  285.85,  285.85,
  285.35,    285.35,  285.35,  285.35,
  284.6,     284.6,   284.6,   284.6,
  284.05,    284.05,  284.05,  284.05,
  283.7,     283.7,   283.7,   283.7,
  283.4,     283.4,   283.4,   283.4,
  283.35,    283.35,  283.35,  283.35,
  283.45,    283.45,  283.45,  283.45,
  283.5,     283.5,   283.5,   283.5,
  283.65,    283.65,  283.65,  283.65,
  283.85,    283.85,  283.85,  283.85,
  284.05,    284.05,  284.05,  284.05,
  284.15,    284.15,  284.15,  284.15,
  284.15,    284.15,  284.15,  284.15,
  284.15,    284.15,  284.15,  284.15,
  284.2,     284.2,   284.2,   284.2,
  284.35,    284.35,  284.35,  284.35,
  284.55,    284.55,  284.55,  284.55,
  284.85,    284.85,  284.85,  284.85,
  285.35,    285.35,  285.35,  285.35,
  286,       286,     286,     286,
  286.6,     286.6,   286.6,   286.6,
  287.05,    287.05,  287.05,  287.05,
  287.45,    287.45,  287.45,  287.45,
  287.85,    287.85,  287.85,  287.85,
  288.2,     288.2,   288.2,   288.2,
  288.5,     288.5,   288.5,   288.5,
  288.6,     288.6,   288.6,   288.6,
  288.75,    288.75,  288.75,  288.75,
  289.05,    289.05,  289.05,  289.05,
  289.15,    289.15,  289.15,  289.15,
  289.15,    289.15,  289.15,  289.15,
  289.1,     289.1,   289.1,   289.1,
  289,       289,     289,     289,
  288.95,    288.95,  288.95,  288.95,
  288.85,    288.85,  288.85,  288.85,
  288.55,    288.55,  288.55,  288.55,
  288.3,     288.3,   288.3,   288.3,
  288.15,    288.15,  288.15,  288.15,
  287.95,    287.95,  287.95,  287.95,
  287.7,     287.7,   287.7,   287.7,
  287.45,    287.45,  287.45,  287.45,
  287.25,    287.25,  287.25,  287.25,
  287,       287,     287,     287,
  286.65,    286.65,  286.65,  286.65,
  286,       286,     286,     286,
  285.2,     285.2,   285.2,   285.2,
  284.45,    284.45,  284.45,  284.45,
  283.8,     283.8,   283.8,   283.8,
  283.45,    283.45,  283.45,  283.45,
  283.2,     283.2,   283.2,   283.2,
  282.95,    282.95,  282.95,  282.95,
  282.8,     282.8,   282.8,   282.8,
  282.8,     282.8,   282.8,   282.8,
  282.9,     282.9,   282.9,   282.9,
  283,       283,     283,     283,
  283.05,    283.05,  283.05,  283.05,
  283,       283,     283,     283,
  282.95,    282.95,  282.95,  282.95,
  283,       283,     283,     283,
  283.05,    283.05,  283.05,  283.05,
  282.95,    282.95,  282.95,  282.95,
  282.85,    282.85,  282.85,  282.85,
  282.7,     282.7,   282.7,   282.7,
  282.5,     282.5,   282.5,   282.5,
  282.85,    282.85,  282.85,  282.85,
  283.9,     283.9,   283.9,   283.9,
  285.15,    285.15,  285.15,  285.15,
  286.3,     286.3,   286.3,   286.3,
  287.7,     287.7,   287.7,   287.7,
  289.2,     289.2,   289.2,   289.2,
  290.3,     290.3,   290.3,   290.3,
  291.1,     291.1,   291.1,   291.1,
  291.65,    291.65,  291.65,  291.65,
  292.05,    292.05,  292.05,  292.05,
  292.45,    292.45,  292.45,  292.45,
  292.7,     292.7,   292.7,   292.7,
  292.75,    292.75,  292.75,  292.75,
  292.9,     292.9,   292.9,   292.9,
  293.15,    293.15,  293.15,  293.15,
  293.3,     293.3,   293.3,   293.3,
  293.35,    293.35,  293.35,  293.35,
  293.4,     293.4,   293.4,   293.4,
  293.3,     293.3,   293.3,   293.3,
  293,       293,     293,     293,
  292.5,     292.5,   292.5,   292.5,
  291.5,     291.5,   291.5,   291.5,
  290.35,    290.35,  290.35,  290.35,
  289.55,    289.55,  289.55,  289.55,
  288.7,     288.7,   288.7,   288.7,
  288.1,     288.1,   288.1,   288.1,
  287.5,     287.5,   287.5,   287.5,
  286.75,    286.75,  286.75,  286.75,
  286.25,    286.25,  286.25,  286.25,
  286.05,    286.05,  286.05,  286.05,
  286.45,    286.45,  286.45,  286.45,
  286.7,     286.7,   286.7,   286.7,
  286.3,     286.3,   286.3,   286.3,
  285.65,    285.65,  285.65,  285.65,
  285.2,     285.2,   285.2,   285.2,
  284.8,     284.8,   284.8,   284.8,
  284.35,    284.35,  284.35,  284.35,
  284,       284,     284,     284,
  283.55,    283.55,  283.55,  283.55,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  283.05,    283.05,  283.05,  283.05,
  282.55,    282.55,  282.55,  282.55,
  282.15,    282.15,  282.15,  282.15,
  282,       282,     282,     282,
  281.8,     281.8,   281.8,   281.8,
  281.65,    281.65,  281.65,  281.65,
  281.8,     281.8,   281.8,   281.8,
  282.45,    282.45,  282.45,  282.45,
  283.6,     283.6,   283.6,   283.6,
  284.6,     284.6,   284.6,   284.6,
  285.35,    285.35,  285.35,  285.35,
  286.1,     286.1,   286.1,   286.1,
  286.9,     286.9,   286.9,   286.9,
  287.9,     287.9,   287.9,   287.9,
  288.85,    288.85,  288.85,  288.85,
  289.75,    289.75,  289.75,  289.75,
  290.8,     290.8,   290.8,   290.8,
  291.7,     291.7,   291.7,   291.7,
  292.3,     292.3,   292.3,   292.3,
  292.65,    292.65,  292.65,  292.65,
  292.95,    292.95,  292.95,  292.95,
  293.25,    293.25,  293.25,  293.25,
  293.4,     293.4,   293.4,   293.4,
  293.45,    293.45,  293.45,  293.45,
  293.3,     293.3,   293.3,   293.3,
  292.9,     292.9,   292.9,   292.9,
  292.35,    292.35,  292.35,  292.35,
  291.7,     291.7,   291.7,   291.7,
  290.95,    290.95,  290.95,  290.95,
  290.15,    290.15,  290.15,  290.15,
  289,       289,     289,     289,
  287.8,     287.8,   287.8,   287.8,
  287.05,    287.05,  287.05,  287.05,
  286.55,    286.55,  286.55,  286.55,
  286.15,    286.15,  286.15,  286.15,
  285.65,    285.65,  285.65,  285.65,
  285.1,     285.1,   285.1,   285.1,
  284.75,    284.75,  284.75,  284.75,
  284.55,    284.55,  284.55,  284.55,
  284.35,    284.35,  284.35,  284.35,
  284.1,     284.1,   284.1,   284.1,
  283.8,     283.8,   283.8,   283.8,
  283.6,     283.6,   283.6,   283.6,
  283.75,    283.75,  283.75,  283.75,
  284.05,    284.05,  284.05,  284.05,
  284.15,    284.15,  284.15,  284.15,
  284.15,    284.15,  284.15,  284.15,
  284.15,    284.15,  284.15,  284.15,
  284.2,     284.2,   284.2,   284.2,
  284.25,    284.25,  284.25,  284.25,
  284.25,    284.25,  284.25,  284.25,
  284.2,     284.2,   284.2,   284.2,
  284.2,     284.2,   284.2,   284.2,
  284.25,    284.25,  284.25,  284.25,
  284.3,     284.3,   284.3,   284.3,
  284.45,    284.45,  284.45,  284.45,
  284.65,    284.65,  284.65,  284.65,
  284.8,     284.8,   284.8,   284.8,
  284.8,     284.8,   284.8,   284.8,
  284.75,    284.75,  284.75,  284.75,
  284.8,     284.8,   284.8,   284.8,
  284.9,     284.9,   284.9,   284.9,
  284.95,    284.95,  284.95,  284.95,
  284.95,    284.95,  284.95,  284.95,
  285.05,    285.05,  285.05,  285.05,
  285.35,    285.35,  285.35,  285.35,
  285.8,     285.8,   285.8,   285.8,
  286.6,     286.6,   286.6,   286.6,
  287.25,    287.25,  287.25,  287.25,
  287.6,     287.6,   287.6,   287.6,
  288,       288,     288,     288,
  288.2,     288.2,   288.2,   288.2,
  288.2,     288.2,   288.2,   288.2,
  288.1,     288.1,   288.1,   288.1,
  287.9,     287.9,   287.9,   287.9,
  287.6,     287.6,   287.6,   287.6,
  287.3,     287.3,   287.3,   287.3,
  286.7,     286.7,   286.7,   286.7,
  285.65,    285.65,  285.65,  285.65,
  284.8,     284.8,   284.8,   284.8,
  284.15,    284.15,  284.15,  284.15,
  283.6,     283.6,   283.6,   283.6,
  283.3,     283.3,   283.3,   283.3,
  282.95,    282.95,  282.95,  282.95,
  282.55,    282.55,  282.55,  282.55,
  282.1,     282.1,   282.1,   282.1,
  281.55,    281.55,  281.55,  281.55,
  280.85,    280.85,  280.85,  280.85,
  280.25,    280.25,  280.25,  280.25,
  280.05,    280.05,  280.05,  280.05,
  279.85,    279.85,  279.85,  279.85,
  279.3,     279.3,   279.3,   279.3,
  278.8,     278.8,   278.8,   278.8,
  278.5,     278.5,   278.5,   278.5,
  278.15,    278.15,  278.15,  278.15,
  277.85,    277.85,  277.85,  277.85,
  277.9,     277.9,   277.9,   277.9,
  278.15,    278.15,  278.15,  278.15,
  278.4,     278.4,   278.4,   278.4,
  278.5,     278.5,   278.5,   278.5,
  278.45,    278.45,  278.45,  278.45,
  278.4,     278.4,   278.4,   278.4,
  278.3,     278.3,   278.3,   278.3,
  278.3,     278.3,   278.3,   278.3,
  278.6,     278.6,   278.6,   278.6,
  279.2,     279.2,   279.2,   279.2,
  279.95,    279.95,  279.95,  279.95,
  280.65,    280.65,  280.65,  280.65,
  281.2,     281.2,   281.2,   281.2,
  281.7,     281.7,   281.7,   281.7,
  282.35,    282.35,  282.35,  282.35,
  283.5,     283.5,   283.5,   283.5,
  285.1,     285.1,   285.1,   285.1,
  287.2,     287.2,   287.2,   287.2,
  288.95,    288.95,  288.95,  288.95,
  289.65,    289.65,  289.65,  289.65,
  290.1,     290.1,   290.1,   290.1,
  290.45,    290.45,  290.45,  290.45,
  290.55,    290.55,  290.55,  290.55,
  290.55,    290.55,  290.55,  290.55,
  290.4,     290.4,   290.4,   290.4,
  289.9,     289.9,   289.9,   289.9,
  289.25,    289.25,  289.25,  289.25,
  288.5,     288.5,   288.5,   288.5,
  287.55,    287.55,  287.55,  287.55,
  286.8,     286.8,   286.8,   286.8,
  286.45,    286.45,  286.45,  286.45,
  286.1,     286.1,   286.1,   286.1,
  285.6,     285.6,   285.6,   285.6,
  285.05,    285.05,  285.05,  285.05,
  284.4,     284.4,   284.4,   284.4,
  283.75,    283.75,  283.75,  283.75,
  282.85,    282.85,  282.85,  282.85,
  282.35,    282.35,  282.35,  282.35,
  282.1,     282.1,   282.1,   282.1,
  280.7,     280.7,   280.7,   280.7,
  279.9,     279.9,   279.9,   279.9,
  279.55,    279.55,  279.55,  279.55,
  278.5,     278.5,   278.5,   278.5,
  277.85,    277.85,  277.85,  277.85,
  277.65,    277.65,  277.65,  277.65,
  277.55,    277.55,  277.55,  277.55,
  277.35,    277.35,  277.35,  277.35,
  277.25,    277.25,  277.25,  277.25,
  277.15,    277.15,  277.15,  277.15,
  277.05,    277.05,  277.05,  277.05,
  277.05,    277.05,  277.05,  277.05,
  277.05,    277.05,  277.05,  277.05,
  277.2,     277.2,   277.2,   277.2,
  277.5,     277.5,   277.5,   277.5,
  277.65,    277.65,  277.65,  277.65,
  277.95,    277.95,  277.95,  277.95,
  278.9,     278.9,   278.9,   278.9,
  280.1,     280.1,   280.1,   280.1,
  281.35,    281.35,  281.35,  281.35,
  282.65,    282.65,  282.65,  282.65,
  283.65,    283.65,  283.65,  283.65,
  284.35,    284.35,  284.35,  284.35,
  285,       285,     285,     285,
  285.9,     285.9,   285.9,   285.9,
  287.15,    287.15,  287.15,  287.15,
  288.2,     288.2,   288.2,   288.2,
  288.75,    288.75,  288.75,  288.75,
  289,       289,     289,     289,
  289.1,     289.1,   289.1,   289.1,
  289.45,    289.45,  289.45,  289.45,
  289.65,    289.65,  289.65,  289.65,
  289.6,     289.6,   289.6,   289.6,
  289.65,    289.65,  289.65,  289.65,
  289.6,     289.6,   289.6,   289.6,
  289.5,     289.5,   289.5,   289.5,
  289.4,     289.4,   289.4,   289.4,
  289.1,     289.1,   289.1,   289.1,
  288.8,     288.8,   288.8,   288.8,
  288.5,     288.5,   288.5,   288.5,
  287.95,    287.95,  287.95,  287.95,
  287.55,    287.55,  287.55,  287.55,
  287.45,    287.45,  287.45,  287.45,
  287.45,    287.45,  287.45,  287.45,
  287.35,    287.35,  287.35,  287.35,
  287.25,    287.25,  287.25,  287.25,
  287.1,     287.1,   287.1,   287.1,
  286.7,     286.7,   286.7,   286.7,
  286.5,     286.5,   286.5,   286.5,
  286.55,    286.55,  286.55,  286.55,
  286.5,     286.5,   286.5,   286.5,
  286.35,    286.35,  286.35,  286.35,
  286.25,    286.25,  286.25,  286.25,
  286.25,    286.25,  286.25,  286.25,
  286.2,     286.2,   286.2,   286.2,
  286.2,     286.2,   286.2,   286.2,
  286.3,     286.3,   286.3,   286.3,
  286.35,    286.35,  286.35,  286.35,
  286.35,    286.35,  286.35,  286.35,
  286.4,     286.4,   286.4,   286.4,
  286.5,     286.5,   286.5,   286.5,
  286.6,     286.6,   286.6,   286.6,
  286.65,    286.65,  286.65,  286.65,
  286.65,    286.65,  286.65,  286.65,
  286.75,    286.75,  286.75,  286.75,
  287,       287,     287,     287,
  287.3,     287.3,   287.3,   287.3,
  287.6,     287.6,   287.6,   287.6,
  287.85,    287.85,  287.85,  287.85,
  288.05,    288.05,  288.05,  288.05,
  288.45,    288.45,  288.45,  288.45,
  289.15,    289.15,  289.15,  289.15,
  289.85,    289.85,  289.85,  289.85,
  290.4,     290.4,   290.4,   290.4,
  290.65,    290.65,  290.65,  290.65,
  290.9,     290.9,   290.9,   290.9,
  291.25,    291.25,  291.25,  291.25,
  291.35,    291.35,  291.35,  291.35,
  291.55,    291.55,  291.55,  291.55,
  291.75,    291.75,  291.75,  291.75,
  291.75,    291.75,  291.75,  291.75,
  291.65,    291.65,  291.65,  291.65,
  291.45,    291.45,  291.45,  291.45,
  291.05,    291.05,  291.05,  291.05,
  290.55,    290.55,  290.55,  290.55,
  290.2,     290.2,   290.2,   290.2,
  289.85,    289.85,  289.85,  289.85,
  289.65,    289.65,  289.65,  289.65,
  289.55,    289.55,  289.55,  289.55,
  289.3,     289.3,   289.3,   289.3,
  289,       289,     289,     289,
  288.45,    288.45,  288.45,  288.45,
  287.7,     287.7,   287.7,   287.7,
  287.2,     287.2,   287.2,   287.2,
  286.95,    286.95,  286.95,  286.95,
  286.75,    286.75,  286.75,  286.75,
  286.6,     286.6,   286.6,   286.6,
  286.55,    286.55,  286.55,  286.55,
  286.6,     286.6,   286.6,   286.6,
  286.65,    286.65,  286.65,  286.65,
  286.65,    286.65,  286.65,  286.65,
  286.7,     286.7,   286.7,   286.7,
  286.75,    286.75,  286.75,  286.75,
  286.75,    286.75,  286.75,  286.75,
  286.75,    286.75,  286.75,  286.75,
  286.8,     286.8,   286.8,   286.8,
  286.85,    286.85,  286.85,  286.85,
  286.9,     286.9,   286.9,   286.9,
  287,       287,     287,     287,
  287.05,    287.05,  287.05,  287.05,
  287.15,    287.15,  287.15,  287.15,
  287.45,    287.45,  287.45,  287.45,
  287.95,    287.95,  287.95,  287.95,
  288.5,     288.5,   288.5,   288.5,
  288.95,    288.95,  288.95,  288.95,
  289.3,     289.3,   289.3,   289.3,
  289.5,     289.5,   289.5,   289.5,
  289.7,     289.7,   289.7,   289.7,
  289.95,    289.95,  289.95,  289.95,
  290.1,     290.1,   290.1,   290.1,
  290.05,    290.05,  290.05,  290.05,
  289.95,    289.95,  289.95,  289.95,
  290.05,    290.05,  290.05,  290.05,
  290.15,    290.15,  290.15,  290.15,
  290.05,    290.05,  290.05,  290.05,
  289.9,     289.9,   289.9,   289.9,
  289.8,     289.8,   289.8,   289.8,
  289.9,     289.9,   289.9,   289.9,
  290.05,    290.05,  290.05,  290.05,
  290,       290,     290,     290,
  289.9,     289.9,   289.9,   289.9,
  289.95,    289.95,  289.95,  289.95,
  290.15,    290.15,  290.15,  290.15,
  290.25,    290.25,  290.25,  290.25,
  290.3,     290.3,   290.3,   290.3,
  290.3,     290.3,   290.3,   290.3,
  290.2,     290.2,   290.2,   290.2,
  290.1,     290.1,   290.1,   290.1,
  290,       290,     290,     290,
  289.9,     289.9,   289.9,   289.9,
  289.7,     289.7,   289.7,   289.7,
  289.4,     289.4,   289.4,   289.4,
  289.15,    289.15,  289.15,  289.15,
  288.8,     288.8,   288.8,   288.8,
  288.45,    288.45,  288.45,  288.45,
  288.25,    288.25,  288.25,  288.25,
  288.1,     288.1,   288.1,   288.1,
  287.95,    287.95,  287.95,  287.95,
  287.75,    287.75,  287.75,  287.75,
  287.55,    287.55,  287.55,  287.55,
  287.35,    287.35,  287.35,  287.35,
  287.15,    287.15,  287.15,  287.15,
  287.05,    287.05,  287.05,  287.05,
  287,       287,     287,     287,
  286.65,    286.65,  286.65,  286.65,
  286.25,    286.25,  286.25,  286.25,
  286.15,    286.15,  286.15,  286.15,
  286.2,     286.2,   286.2,   286.2,
  286.3,     286.3,   286.3,   286.3,
  286.4,     286.4,   286.4,   286.4,
  286.45,    286.45,  286.45,  286.45,
  286.5,     286.5,   286.5,   286.5,
  286.75,    286.75,  286.75,  286.75,
  286.95,    286.95,  286.95,  286.95,
  286.95,    286.95,  286.95,  286.95,
  287,       287,     287,     287,
  286.6,     286.6,   286.6,   286.6,
  286.45,    286.45,  286.45,  286.45,
  286.55,    286.55,  286.55,  286.55,
  286.3,     286.3,   286.3,   286.3,
  287.1,     287.1,   287.1,   287.1,
  287.75,    287.75,  287.75,  287.75,
  287.6,     287.6,   287.6,   287.6,
  287.95,    287.95,  287.95,  287.95,
  287.85,    287.85,  287.85,  287.85,
  287.1,     287.1,   287.1,   287.1,
  286.55,    286.55,  286.55,  286.55,
  285.9,     285.9,   285.9,   285.9,
  285.2,     285.2,   285.2,   285.2,
  284.75,    284.75,  284.75,  284.75,
  284.4,     284.4,   284.4,   284.4,
  284.45,    284.45,  284.45,  284.45,
  284.7,     284.7,   284.7,   284.7,
  284.5,     284.5,   284.5,   284.5,
  284.1,     284.1,   284.1,   284.1,
  283.85,    283.85,  283.85,  283.85,
  283.7,     283.7,   283.7,   283.7,
  283.55,    283.55,  283.55,  283.55,
  283.35,    283.35,  283.35,  283.35,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.2,     283.2,   283.2,   283.2,
  283.05,    283.05,  283.05,  283.05,
  282.85,    282.85,  282.85,  282.85,
  282.6,     282.6,   282.6,   282.6,
  282.05,    282.05,  282.05,  282.05,
  281.45,    281.45,  281.45,  281.45,
  281,       281,     281,     281,
  280.7,     280.7,   280.7,   280.7,
  280.55,    280.55,  280.55,  280.55,
  280.5,     280.5,   280.5,   280.5,
  280.45,    280.45,  280.45,  280.45,
  280.2,     280.2,   280.2,   280.2,
  279.9,     279.9,   279.9,   279.9,
  279.55,    279.55,  279.55,  279.55,
  279.45,    279.45,  279.45,  279.45,
  279.55,    279.55,  279.55,  279.55,
  279.55,    279.55,  279.55,  279.55,
  279.55,    279.55,  279.55,  279.55,
  279.8,     279.8,   279.8,   279.8,
  280.65,    280.65,  280.65,  280.65,
  282.3,     282.3,   282.3,   282.3,
  283.95,    283.95,  283.95,  283.95,
  284.95,    284.95,  284.95,  284.95,
  285.85,    285.85,  285.85,  285.85,
  286.45,    286.45,  286.45,  286.45,
  286.8,     286.8,   286.8,   286.8,
  287.1,     287.1,   287.1,   287.1,
  286.9,     286.9,   286.9,   286.9,
  286.85,    286.85,  286.85,  286.85,
  287.4,     287.4,   287.4,   287.4,
  287.75,    287.75,  287.75,  287.75,
  287.55,    287.55,  287.55,  287.55,
  287.45,    287.45,  287.45,  287.45,
  287.6,     287.6,   287.6,   287.6,
  287.45,    287.45,  287.45,  287.45,
  287.15,    287.15,  287.15,  287.15,
  287.05,    287.05,  287.05,  287.05,
  286.8,     286.8,   286.8,   286.8,
  286.4,     286.4,   286.4,   286.4,
  286.3,     286.3,   286.3,   286.3,
  286.3,     286.3,   286.3,   286.3,
  286.1,     286.1,   286.1,   286.1,
  285.95,    285.95,  285.95,  285.95,
  285.75,    285.75,  285.75,  285.75,
  285.25,    285.25,  285.25,  285.25,
  284.75,    284.75,  284.75,  284.75,
  284.65,    284.65,  284.65,  284.65,
  284.95,    284.95,  284.95,  284.95,
  285.3,     285.3,   285.3,   285.3,
  285.5,     285.5,   285.5,   285.5,
  285.65,    285.65,  285.65,  285.65,
  285.7,     285.7,   285.7,   285.7,
  285.65,    285.65,  285.65,  285.65,
  285.65,    285.65,  285.65,  285.65,
  285.7,     285.7,   285.7,   285.7,
  285.75,    285.75,  285.75,  285.75,
  285.85,    285.85,  285.85,  285.85,
  286,       286,     286,     286,
  286,       286,     286,     286,
  285.95,    285.95,  285.95,  285.95,
  285.95,    285.95,  285.95,  285.95,
  286.05,    286.05,  286.05,  286.05,
  286.2,     286.2,   286.2,   286.2,
  286.2,     286.2,   286.2,   286.2,
  286.1,     286.1,   286.1,   286.1,
  286.05,    286.05,  286.05,  286.05,
  286.15,    286.15,  286.15,  286.15,
  286.3,     286.3,   286.3,   286.3,
  286.6,     286.6,   286.6,   286.6,
  287.3,     287.3,   287.3,   287.3,
  287.85,    287.85,  287.85,  287.85,
  288.5,     288.5,   288.5,   288.5,
  289.1,     289.1,   289.1,   289.1,
  289.2,     289.2,   289.2,   289.2,
  289.3,     289.3,   289.3,   289.3,
  289.4,     289.4,   289.4,   289.4,
  289.5,     289.5,   289.5,   289.5,
  289.45,    289.45,  289.45,  289.45,
  289.35,    289.35,  289.35,  289.35,
  289.3,     289.3,   289.3,   289.3,
  289.25,    289.25,  289.25,  289.25,
  289.2,     289.2,   289.2,   289.2,
  289.05,    289.05,  289.05,  289.05,
  288.95,    288.95,  288.95,  288.95,
  288.9,     288.9,   288.9,   288.9,
  288.8,     288.8,   288.8,   288.8,
  288.7,     288.7,   288.7,   288.7,
  288.45,    288.45,  288.45,  288.45,
  288.2,     288.2,   288.2,   288.2,
  287.9,     287.9,   287.9,   287.9,
  287.35,    287.35,  287.35,  287.35,
  286.9,     286.9,   286.9,   286.9,
  286.55,    286.55,  286.55,  286.55,
  286.25,    286.25,  286.25,  286.25,
  286,       286,     286,     286,
  285.7,     285.7,   285.7,   285.7,
  285.6,     285.6,   285.6,   285.6,
  285.65,    285.65,  285.65,  285.65,
  285.6,     285.6,   285.6,   285.6,
  285.5,     285.5,   285.5,   285.5,
  285.35,    285.35,  285.35,  285.35,
  285.2,     285.2,   285.2,   285.2,
  285.1,     285.1,   285.1,   285.1,
  285.05,    285.05,  285.05,  285.05,
  285.05,    285.05,  285.05,  285.05,
  285.2,     285.2,   285.2,   285.2,
  285.5,     285.5,   285.5,   285.5,
  285.7,     285.7,   285.7,   285.7,
  285.7,     285.7,   285.7,   285.7,
  285.6,     285.6,   285.6,   285.6,
  285.55,    285.55,  285.55,  285.55,
  285.65,    285.65,  285.65,  285.65,
  285.7,     285.7,   285.7,   285.7,
  285.6,     285.6,   285.6,   285.6,
  285.55,    285.55,  285.55,  285.55,
  285.5,     285.5,   285.5,   285.5,
  285.45,    285.45,  285.45,  285.45,
  285.55,    285.55,  285.55,  285.55,
  285.65,    285.65,  285.65,  285.65,
  285.7,     285.7,   285.7,   285.7,
  285.9,     285.9,   285.9,   285.9,
  286.2,     286.2,   286.2,   286.2,
  286.7,     286.7,   286.7,   286.7,
  287.4,     287.4,   287.4,   287.4,
  288.1,     288.1,   288.1,   288.1,
  288.7,     288.7,   288.7,   288.7,
  288.95,    288.95,  288.95,  288.95,
  288.9,     288.9,   288.9,   288.9,
  288.85,    288.85,  288.85,  288.85,
  288.85,    288.85,  288.85,  288.85,
  288.75,    288.75,  288.75,  288.75,
  288.55,    288.55,  288.55,  288.55,
  288.25,    288.25,  288.25,  288.25,
  287.95,    287.95,  287.95,  287.95,
  287.7,     287.7,   287.7,   287.7,
  287.45,    287.45,  287.45,  287.45,
  287.3,     287.3,   287.3,   287.3,
  287.2,     287.2,   287.2,   287.2,
  287.05,    287.05,  287.05,  287.05,
  286.85,    286.85,  286.85,  286.85,
  286.7,     286.7,   286.7,   286.7,
  286.6,     286.6,   286.6,   286.6,
  286.5,     286.5,   286.5,   286.5,
  286.45,    286.45,  286.45,  286.45,
  286.45,    286.45,  286.45,  286.45,
  286.4,     286.4,   286.4,   286.4,
  286.35,    286.35,  286.35,  286.35,
  286.3,     286.3,   286.3,   286.3,
  286.25,    286.25,  286.25,  286.25,
  286.15,    286.15,  286.15,  286.15,
  286.05,    286.05,  286.05,  286.05,
  285.95,    285.95,  285.95,  285.95,
  285.7,     285.7,   285.7,   285.7,
  285.35,    285.35,  285.35,  285.35,
  284.8,     284.8,   284.8,   284.8,
  284.1,     284.1,   284.1,   284.1,
  283.45,    283.45,  283.45,  283.45,
  282.95,    282.95,  282.95,  282.95,
  282.7,     282.7,   282.7,   282.7,
  282.6,     282.6,   282.6,   282.6,
  282.5,     282.5,   282.5,   282.5,
  282.6,     282.6,   282.6,   282.6,
  283.1,     283.1,   283.1,   283.1,
  283.85,    283.85,  283.85,  283.85,
  284.8,     284.8,   284.8,   284.8,
  286.05,    286.05,  286.05,  286.05,
  287.05,    287.05,  287.05,  287.05,
  287.9,     287.9,   287.9,   287.9,
  289,       289,     289,     289,
  290,       290,     290,     290,
  290.65,    290.65,  290.65,  290.65,
  291,       291,     291,     291,
  291.35,    291.35,  291.35,  291.35,
  291.85,    291.85,  291.85,  291.85,
  292.4,     292.4,   292.4,   292.4,
  292.5,     292.5,   292.5,   292.5,
  292.45,    292.45,  292.45,  292.45,
  292.7,     292.7,   292.7,   292.7,
  292.95,    292.95,  292.95,  292.95,
  292.8,     292.8,   292.8,   292.8,
  292.3,     292.3,   292.3,   292.3,
  291.7,     291.7,   291.7,   291.7,
  291.15,    291.15,  291.15,  291.15,
  290.9,     290.9,   290.9,   290.9,
  290.9,     290.9,   290.9,   290.9,
  290.9,     290.9,   290.9,   290.9,
  290.8,     290.8,   290.8,   290.8,
  290.6,     290.6,   290.6,   290.6,
  290.25,    290.25,  290.25,  290.25,
  289.95,    289.95,  289.95,  289.95,
  289.7,     289.7,   289.7,   289.7,
  289.45,    289.45,  289.45,  289.45,
  289.4,     289.4,   289.4,   289.4,
  289.55,    289.55,  289.55,  289.55,
  289.8,     289.8,   289.8,   289.8,
  290.15,    290.15,  290.15,  290.15,
  290.4,     290.4,   290.4,   290.4,
  290.4,     290.4,   290.4,   290.4,
  289.85,    289.85,  289.85,  289.85,
  289.25,    289.25,  289.25,  289.25,
  289.05,    289.05,  289.05,  289.05,
  288.9,     288.9,   288.9,   288.9,
  288.8,     288.8,   288.8,   288.8,
  288.75,    288.75,  288.75,  288.75,
  288.8,     288.8,   288.8,   288.8,
  288.85,    288.85,  288.85,  288.85,
  288.85,    288.85,  288.85,  288.85,
  288.9,     288.9,   288.9,   288.9,
  289,       289,     289,     289,
  289.05,    289.05,  289.05,  289.05,
  289.1,     289.1,   289.1,   289.1,
  289.15,    289.15,  289.15,  289.15,
  289.2,     289.2,   289.2,   289.2,
  289.4,     289.4,   289.4,   289.4,
  289.75,    289.75,  289.75,  289.75,
  290.15,    290.15,  290.15,  290.15,
  290.55,    290.55,  290.55,  290.55,
  291.2,     291.2,   291.2,   291.2,
  291.95,    291.95,  291.95,  291.95,
  292.4,     292.4,   292.4,   292.4,
  292.7,     292.7,   292.7,   292.7,
  290.75,    290.75,  290.75,  290.75,
  287.85,    287.85,  287.85,  287.85,
  288.05,    288.05,  288.05,  288.05,
  289.1,     289.1,   289.1,   289.1,
  287.6,     287.6,   287.6,   287.6,
  285.9,     285.9,   285.9,   285.9,
  286,       286,     286,     286,
  286.3,     286.3,   286.3,   286.3,
  286.3,     286.3,   286.3,   286.3,
  286.2,     286.2,   286.2,   286.2,
  286.15,    286.15,  286.15,  286.15,
  286.2,     286.2,   286.2,   286.2,
  286.35,    286.35,  286.35,  286.35,
  286.3,     286.3,   286.3,   286.3,
  286.2,     286.2,   286.2,   286.2,
  286.1,     286.1,   286.1,   286.1,
  285.85,    285.85,  285.85,  285.85,
  285.8,     285.8,   285.8,   285.8,
  285.75,    285.75,  285.75,  285.75,
  285.55,    285.55,  285.55,  285.55,
  285.4,     285.4,   285.4,   285.4,
  285.5,     285.5,   285.5,   285.5,
  285.65,    285.65,  285.65,  285.65,
  285.5,     285.5,   285.5,   285.5,
  285.2,     285.2,   285.2,   285.2,
  285.15,    285.15,  285.15,  285.15,
  285.2,     285.2,   285.2,   285.2,
  285.15,    285.15,  285.15,  285.15,
  285.3,     285.3,   285.3,   285.3,
  285.6,     285.6,   285.6,   285.6,
  285.8,     285.8,   285.8,   285.8,
  285.8,     285.8,   285.8,   285.8,
  285.85,    285.85,  285.85,  285.85,
  286,       286,     286,     286,
  286.05,    286.05,  286.05,  286.05,
  286,       286,     286,     286,
  286.05,    286.05,  286.05,  286.05,
  286.4,     286.4,   286.4,   286.4,
  286.7,     286.7,   286.7,   286.7,
  286.4,     286.4,   286.4,   286.4,
  285.65,    285.65,  285.65,  285.65,
  285.5,     285.5,   285.5,   285.5,
  286,       286,     286,     286,
  286.55,    286.55,  286.55,  286.55,
  287.15,    287.15,  287.15,  287.15,
  287.65,    287.65,  287.65,  287.65,
  288.05,    288.05,  288.05,  288.05,
  288.35,    288.35,  288.35,  288.35,
  288.6,     288.6,   288.6,   288.6,
  288.95,    288.95,  288.95,  288.95,
  289.15,    289.15,  289.15,  289.15,
  289.3,     289.3,   289.3,   289.3,
  289.55,    289.55,  289.55,  289.55,
  289.65,    289.65,  289.65,  289.65,
  289.35,    289.35,  289.35,  289.35,
  288.9,     288.9,   288.9,   288.9,
  288.75,    288.75,  288.75,  288.75,
  288.6,     288.6,   288.6,   288.6,
  288.25,    288.25,  288.25,  288.25,
  288.05,    288.05,  288.05,  288.05,
  288.15,    288.15,  288.15,  288.15,
  288.35,    288.35,  288.35,  288.35,
  288.5,     288.5,   288.5,   288.5,
  288.65,    288.65,  288.65,  288.65,
  288.95,    288.95,  288.95,  288.95,
  289.3,     289.3,   289.3,   289.3,
  289.65,    289.65,  289.65,  289.65,
  290,       290,     290,     290,
  290.3,     290.3,   290.3,   290.3,
  290.55,    290.55,  290.55,  290.55,
  290.65,    290.65,  290.65,  290.65,
  290.65,    290.65,  290.65,  290.65,
  290.6,     290.6,   290.6,   290.6,
  290.5,     290.5,   290.5,   290.5,
  290.3,     290.3,   290.3,   290.3,
  290.15,    290.15,  290.15,  290.15,
  290.1,     290.1,   290.1,   290.1,
  290.05,    290.05,  290.05,  290.05,
  290.15,    290.15,  290.15,  290.15,
  290.2,     290.2,   290.2,   290.2,
  290.05,    290.05,  290.05,  290.05,
  289.95,    289.95,  289.95,  289.95,
  289.95,    289.95,  289.95,  289.95,
  290.05,    290.05,  290.05,  290.05,
  290.25,    290.25,  290.25,  290.25,
  290.55,    290.55,  290.55,  290.55,
  290.9,     290.9,   290.9,   290.9,
  290.95,    290.95,  290.95,  290.95,
  290.95,    290.95,  290.95,  290.95,
  291.05,    291.05,  291.05,  291.05,
  291.05,    291.05,  291.05,  291.05,
  290.9,     290.9,   290.9,   290.9,
  290.85,    290.85,  290.85,  290.85,
  291.05,    291.05,  291.05,  291.05,
  290.5,     290.5,   290.5,   290.5,
  289.75,    289.75,  289.75,  289.75,
  290.2,     290.2,   290.2,   290.2,
  290.9,     290.9,   290.9,   290.9,
  291,       291,     291,     291,
  290.9,     290.9,   290.9,   290.9,
  290.8,     290.8,   290.8,   290.8,
  290.65,    290.65,  290.65,  290.65,
  290.5,     290.5,   290.5,   290.5,
  290.35,    290.35,  290.35,  290.35,
  290.2,     290.2,   290.2,   290.2,
  290.2,     290.2,   290.2,   290.2,
  290.15,    290.15,  290.15,  290.15,
  289.85,    289.85,  289.85,  289.85,
  289.45,    289.45,  289.45,  289.45,
  289.15,    289.15,  289.15,  289.15,
  288.9,     288.9,   288.9,   288.9,
  288.65,    288.65,  288.65,  288.65,
  288.45,    288.45,  288.45,  288.45,
  288.3,     288.3,   288.3,   288.3,
  288.35,    288.35,  288.35,  288.35,
  288.5,     288.5,   288.5,   288.5,
  288.65,    288.65,  288.65,  288.65,
  288.85,    288.85,  288.85,  288.85,
  288.7,     288.7,   288.7,   288.7,
  288.45,    288.45,  288.45,  288.45,
  288.5,     288.5,   288.5,   288.5,
  288.55,    288.55,  288.55,  288.55,
  288.45,    288.45,  288.45,  288.45,
  288.35,    288.35,  288.35,  288.35,
  288.3,     288.3,   288.3,   288.3,
  288.25,    288.25,  288.25,  288.25,
  288.1,     288.1,   288.1,   288.1,
  287.95,    287.95,  287.95,  287.95,
  287.8,     287.8,   287.8,   287.8,
  287.6,     287.6,   287.6,   287.6,
  287.65,    287.65,  287.65,  287.65,
  287.75,    287.75,  287.75,  287.75,
  287.75,    287.75,  287.75,  287.75,
  287.8,     287.8,   287.8,   287.8,
  287.8,     287.8,   287.8,   287.8,
  287.4,     287.4,   287.4,   287.4,
  287.05,    287.05,  287.05,  287.05,
  287.2,     287.2,   287.2,   287.2,
  287.3,     287.3,   287.3,   287.3,
  287.25,    287.25,  287.25,  287.25,
  287.25,    287.25,  287.25,  287.25,
  287.4,     287.4,   287.4,   287.4,
  287.45,    287.45,  287.45,  287.45,
  287.3,     287.3,   287.3,   287.3,
  287.35,    287.35,  287.35,  287.35,
  287.75,    287.75,  287.75,  287.75,
  287.85,    287.85,  287.85,  287.85,
  287.55,    287.55,  287.55,  287.55,
  287.45,    287.45,  287.45,  287.45,
  287.4,     287.4,   287.4,   287.4,
  287.15,    287.15,  287.15,  287.15,
  286.95,    286.95,  286.95,  286.95,
  286.75,    286.75,  286.75,  286.75,
  285.85,    285.85,  285.85,  285.85,
  285,       285,     285,     285,
  284.7,     284.7,   284.7,   284.7,
  284.4,     284.4,   284.4,   284.4,
  284.25,    284.25,  284.25,  284.25,
  284.15,    284.15,  284.15,  284.15,
  284.2,     284.2,   284.2,   284.2,
  284.05,    284.05,  284.05,  284.05,
  283.7,     283.7,   283.7,   283.7,
  283.6,     283.6,   283.6,   283.6,
  283.7,     283.7,   283.7,   283.7,
  283.85,    283.85,  283.85,  283.85,
  283.85,    283.85,  283.85,  283.85,
  283.75,    283.75,  283.75,  283.75,
  283.7,     283.7,   283.7,   283.7,
  283.7,     283.7,   283.7,   283.7,
  283.6,     283.6,   283.6,   283.6,
  283.6,     283.6,   283.6,   283.6,
  283.9,     283.9,   283.9,   283.9,
  284.2,     284.2,   284.2,   284.2,
  284.25,    284.25,  284.25,  284.25,
  284.25,    284.25,  284.25,  284.25,
  284.25,    284.25,  284.25,  284.25,
  284.25,    284.25,  284.25,  284.25,
  284.15,    284.15,  284.15,  284.15,
  284.05,    284.05,  284.05,  284.05,
  284.15,    284.15,  284.15,  284.15,
  284.3,     284.3,   284.3,   284.3,
  284.25,    284.25,  284.25,  284.25,
  283.85,    283.85,  283.85,  283.85,
  283.55,    283.55,  283.55,  283.55,
  283.65,    283.65,  283.65,  283.65,
  283.85,    283.85,  283.85,  283.85,
  284.1,     284.1,   284.1,   284.1,
  285.05,    285.05,  285.05,  285.05,
  286,       286,     286,     286,
  286.35,    286.35,  286.35,  286.35,
  286.4,     286.4,   286.4,   286.4,
  286.5,     286.5,   286.5,   286.5,
  286.85,    286.85,  286.85,  286.85,
  286.85,    286.85,  286.85,  286.85,
  286.45,    286.45,  286.45,  286.45,
  285.25,    285.25,  285.25,  285.25,
  284.65,    284.65,  284.65,  284.65,
  285,       285,     285,     285,
  285.05,    285.05,  285.05,  285.05,
  285,       285,     285,     285,
  284.8,     284.8,   284.8,   284.8,
  284.45,    284.45,  284.45,  284.45,
  284.05,    284.05,  284.05,  284.05,
  283.7,     283.7,   283.7,   283.7,
  283.45,    283.45,  283.45,  283.45,
  283.3,     283.3,   283.3,   283.3,
  283.15,    283.15,  283.15,  283.15,
  283,       283,     283,     283,
  282.85,    282.85,  282.85,  282.85,
  282.65,    282.65,  282.65,  282.65,
  282.45,    282.45,  282.45,  282.45,
  282.3,     282.3,   282.3,   282.3,
  282.25,    282.25,  282.25,  282.25,
  282.2,     282.2,   282.2,   282.2,
  282.15,    282.15,  282.15,  282.15,
  282.15,    282.15,  282.15,  282.15,
  282.1,     282.1,   282.1,   282.1,
  281.95,    281.95,  281.95,  281.95,
  281.6,     281.6,   281.6,   281.6,
  281.1,     281.1,   281.1,   281.1,
  280.5,     280.5,   280.5,   280.5,
  279.95,    279.95,  279.95,  279.95,
  279.7,     279.7,   279.7,   279.7,
  279.45,    279.45,  279.45,  279.45,
  279.1,     279.1,   279.1,   279.1,
  279.05,    279.05,  279.05,  279.05,
  279,       279,     279,     279,
  278.8,     278.8,   278.8,   278.8,
  278.85,    278.85,  278.85,  278.85,
  279.65,    279.65,  279.65,  279.65,
  281.2,     281.2,   281.2,   281.2,
  282.65,    282.65,  282.65,  282.65,
  283.9,     283.9,   283.9,   283.9,
  284.9,     284.9,   284.9,   284.9,
  284.8,     284.8,   284.8,   284.8,
  284.4,     284.4,   284.4,   284.4,
  284.15,    284.15,  284.15,  284.15,
  283.65,    283.65,  283.65,  283.65,
  284.1,     284.1,   284.1,   284.1,
  284.9,     284.9,   284.9,   284.9,
  285.25,    285.25,  285.25,  285.25,
  285.15,    285.15,  285.15,  285.15,
  284.2,     284.2,   284.2,   284.2,
  283,       283,     283,     283,
  283.1,     283.1,   283.1,   283.1,
  283.9,     283.9,   283.9,   283.9,
  283.9,     283.9,   283.9,   283.9,
  283.7,     283.7,   283.7,   283.7,
  283.2,     283.2,   283.2,   283.2,
  282.25,    282.25,  282.25,  282.25,
  281.45,    281.45,  281.45,  281.45,
  281.05,    281.05,  281.05,  281.05,
  281,       281,     281,     281,
  281.1,     281.1,   281.1,   281.1,
  281.3,     281.3,   281.3,   281.3,
  281.35,    281.35,  281.35,  281.35,
  281.05,    281.05,  281.05,  281.05,
  280.65,    280.65,  280.65,  280.65,
  280.3,     280.3,   280.3,   280.3,
  280,       280,     280,     280,
  279.75,    279.75,  279.75,  279.75,
  279.55,    279.55,  279.55,  279.55,
  279.35,    279.35,  279.35,  279.35,
  279.15,    279.15,  279.15,  279.15,
  279.2,     279.2,   279.2,   279.2,
  279.45,    279.45,  279.45,  279.45,
  279.8,     279.8,   279.8,   279.8,
  280.25,    280.25,  280.25,  280.25,
  280.55,    280.55,  280.55,  280.55,
  280.5,     280.5,   280.5,   280.5,
  280.25,    280.25,  280.25,  280.25,
  280.15,    280.15,  280.15,  280.15,
  280.15,    280.15,  280.15,  280.15,
  280.15,    280.15,  280.15,  280.15,
  280.15,    280.15,  280.15,  280.15,
  280.15,    280.15,  280.15,  280.15,
  280.15,    280.15,  280.15,  280.15,
  280.2,     280.2,   280.2,   280.2,
  280.55,    280.55,  280.55,  280.55,
  281.15,    281.15,  281.15,  281.15,
  281.65,    281.65,  281.65,  281.65,
  282.2,     282.2,   282.2,   282.2,
  281.25,    281.25,  281.25,  281.25,
  279.8,     279.8,   279.8,   279.8,
  279.9,     279.9,   279.9,   279.9,
  280.4,     280.4,   280.4,   280.4,
  280.85,    280.85,  280.85,  280.85,
  281.75,    281.75,  281.75,  281.75,
  282.45,    282.45,  282.45,  282.45,
  282.1,     282.1,   282.1,   282.1,
  282.05,    282.05,  282.05,  282.05,
  282.4,     282.4,   282.4,   282.4,
  282.55,    282.55,  282.55,  282.55,
  282.55,    282.55,  282.55,  282.55,
  282.25,    282.25,  282.25,  282.25,
  281.95,    281.95,  281.95,  281.95,
  281.6,     281.6,   281.6,   281.6,
  281.1,     281.1,   281.1,   281.1,
  280.85,    280.85,  280.85,  280.85,
  280.9,     280.9,   280.9,   280.9,
  281,       281,     281,     281,
  281.05,    281.05,  281.05,  281.05,
  281,       281,     281,     281,
  280.85,    280.85,  280.85,  280.85,
  280.7,     280.7,   280.7,   280.7,
  280.7,     280.7,   280.7,   280.7,
  280.8,     280.8,   280.8,   280.8,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.6,     280.6,   280.6,   280.6,
  280.65,    280.65,  280.65,  280.65,
  280.65,    280.65,  280.65,  280.65,
  280.45,    280.45,  280.45,  280.45,
  280.4,     280.4,   280.4,   280.4,
  280.3,     280.3,   280.3,   280.3,
  279.9,     279.9,   279.9,   279.9,
  279.7,     279.7,   279.7,   279.7,
  279.8,     279.8,   279.8,   279.8,
  279.65,    279.65,  279.65,  279.65,
  279.25,    279.25,  279.25,  279.25,
  279.1,     279.1,   279.1,   279.1,
  279.05,    279.05,  279.05,  279.05,
  279.2,     279.2,   279.2,   279.2,
  279.85,    279.85,  279.85,  279.85,
  280.45,    280.45,  280.45,  280.45,
  280.9,     280.9,   280.9,   280.9,
  281.75,    281.75,  281.75,  281.75,
  282.55,    282.55,  282.55,  282.55,
  282.9,     282.9,   282.9,   282.9,
  283.2,     283.2,   283.2,   283.2,
  283.6,     283.6,   283.6,   283.6,
  284.05,    284.05,  284.05,  284.05,
  284.3,     284.3,   284.3,   284.3,
  284.25,    284.25,  284.25,  284.25,
  283.9,     283.9,   283.9,   283.9,
  282.95,    282.95,  282.95,  282.95,
  282.35,    282.35,  282.35,  282.35,
  282.65,    282.65,  282.65,  282.65,
  282.75,    282.75,  282.75,  282.75,
  282.6,     282.6,   282.6,   282.6,
  282.5,     282.5,   282.5,   282.5,
  282.3,     282.3,   282.3,   282.3,
  282,       282,     282,     282,
  281.7,     281.7,   281.7,   281.7,
  281.35,    281.35,  281.35,  281.35,
  281.05,    281.05,  281.05,  281.05,
  280.9,     280.9,   280.9,   280.9,
  280.85,    280.85,  280.85,  280.85,
  280.85,    280.85,  280.85,  280.85,
  280.8,     280.8,   280.8,   280.8,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.6,     280.6,   280.6,   280.6,
  280.55,    280.55,  280.55,  280.55,
  280.6,     280.6,   280.6,   280.6,
  280.6,     280.6,   280.6,   280.6,
  280.55,    280.55,  280.55,  280.55,
  280.5,     280.5,   280.5,   280.5,
  280.45,    280.45,  280.45,  280.45,
  280.45,    280.45,  280.45,  280.45,
  280.4,     280.4,   280.4,   280.4,
  280.35,    280.35,  280.35,  280.35,
  280.35,    280.35,  280.35,  280.35,
  280.35,    280.35,  280.35,  280.35,
  280.35,    280.35,  280.35,  280.35,
  280.35,    280.35,  280.35,  280.35,
  280.3,     280.3,   280.3,   280.3,
  280.2,     280.2,   280.2,   280.2,
  280.05,    280.05,  280.05,  280.05,
  279.9,     279.9,   279.9,   279.9,
  279.8,     279.8,   279.8,   279.8,
  279.7,     279.7,   279.7,   279.7,
  279.7,     279.7,   279.7,   279.7,
  279.8,     279.8,   279.8,   279.8,
  279.95,    279.95,  279.95,  279.95,
  280.1,     280.1,   280.1,   280.1,
  280.15,    280.15,  280.15,  280.15,
  280.35,    280.35,  280.35,  280.35,
  280.55,    280.55,  280.55,  280.55,
  280.7,     280.7,   280.7,   280.7,
  281,       281,     281,     281,
  281.3,     281.3,   281.3,   281.3,
  281.65,    281.65,  281.65,  281.65,
  281.9,     281.9,   281.9,   281.9,
  282,       282,     282,     282,
  282.3,     282.3,   282.3,   282.3,
  282.55,    282.55,  282.55,  282.55,
  282.45,    282.45,  282.45,  282.45,
  282.25,    282.25,  282.25,  282.25,
  282,       282,     282,     282,
  281.7,     281.7,   281.7,   281.7,
  281.45,    281.45,  281.45,  281.45,
  281.3,     281.3,   281.3,   281.3,
  280.9,     280.9,   280.9,   280.9,
  280.15,    280.15,  280.15,  280.15,
  279.6,     279.6,   279.6,   279.6,
  279.4,     279.4,   279.4,   279.4,
  279.5,     279.5,   279.5,   279.5,
  279.3,     279.3,   279.3,   279.3,
  278.8,     278.8,   278.8,   278.8,
  278.8,     278.8,   278.8,   278.8,
  279.2,     279.2,   279.2,   279.2,
  279.3,     279.3,   279.3,   279.3,
  279.4,     279.4,   279.4,   279.4,
  279.45,    279.45,  279.45,  279.45,
  279.25,    279.25,  279.25,  279.25,
  279.1,     279.1,   279.1,   279.1,
  278.85,    278.85,  278.85,  278.85,
  278.7,     278.7,   278.7,   278.7,
  278.55,    278.55,  278.55,  278.55,
  278.25,    278.25,  278.25,  278.25,
  277.9,     277.9,   277.9,   277.9,
  277.7,     277.7,   277.7,   277.7,
  277.6,     277.6,   277.6,   277.6,
  277.6,     277.6,   277.6,   277.6,
  277.75,    277.75,  277.75,  277.75,
  277.9,     277.9,   277.9,   277.9,
  278.05,    278.05,  278.05,  278.05,
  278.2,     278.2,   278.2,   278.2,
  278.35,    278.35,  278.35,  278.35,
  278.65,    278.65,  278.65,  278.65,
  278.95,    278.95,  278.95,  278.95,
  279.25,    279.25,  279.25,  279.25,
  279.5,     279.5,   279.5,   279.5,
  279.55,    279.55,  279.55,  279.55,
  279.75,    279.75,  279.75,  279.75,
  280.35,    280.35,  280.35,  280.35,
  280.95,    280.95,  280.95,  280.95,
  281.25,    281.25,  281.25,  281.25,
  281.5,     281.5,   281.5,   281.5,
  281.85,    281.85,  281.85,  281.85,
  282.25,    282.25,  282.25,  282.25,
  282.55,    282.55,  282.55,  282.55,
  282.75,    282.75,  282.75,  282.75,
  282.95,    282.95,  282.95,  282.95,
  283.05,    283.05,  283.05,  283.05,
  282.9,     282.9,   282.9,   282.9,
  282.6,     282.6,   282.6,   282.6,
  282.25,    282.25,  282.25,  282.25,
  281.85,    281.85,  281.85,  281.85,
  281.55,    281.55,  281.55,  281.55,
  281.3,     281.3,   281.3,   281.3,
  281.1,     281.1,   281.1,   281.1,
  280.95,    280.95,  280.95,  280.95,
  280.8,     280.8,   280.8,   280.8,
  280.8,     280.8,   280.8,   280.8,
  280.85,    280.85,  280.85,  280.85,
  280.85,    280.85,  280.85,  280.85,
  280.8,     280.8,   280.8,   280.8,
  280.85,    280.85,  280.85,  280.85,
  281,       281,     281,     281,
  281.15,    281.15,  281.15,  281.15,
  281.35,    281.35,  281.35,  281.35,
  281.5,     281.5,   281.5,   281.5,
  281.6,     281.6,   281.6,   281.6,
  281.75,    281.75,  281.75,  281.75,
  281.9,     281.9,   281.9,   281.9,
  282,       282,     282,     282,
  282.15,    282.15,  282.15,  282.15,
  282.3,     282.3,   282.3,   282.3,
  282.4,     282.4,   282.4,   282.4,
  282.45,    282.45,  282.45,  282.45,
  282.6,     282.6,   282.6,   282.6,
  282.75,    282.75,  282.75,  282.75,
  282.75,    282.75,  282.75,  282.75,
  282.75,    282.75,  282.75,  282.75,
  282.85,    282.85,  282.85,  282.85,
  283.05,    283.05,  283.05,  283.05,
  283.25,    283.25,  283.25,  283.25,
  283.45,    283.45,  283.45,  283.45,
  283.7,     283.7,   283.7,   283.7,
  284.1,     284.1,   284.1,   284.1,
  284.65,    284.65,  284.65,  284.65,
  285.3,     285.3,   285.3,   285.3,
  285.95,    285.95,  285.95,  285.95,
  286.55,    286.55,  286.55,  286.55,
  287.2,     287.2,   287.2,   287.2,
  287.85,    287.85,  287.85,  287.85,
  288.4,     288.4,   288.4,   288.4,
  288.65,    288.65,  288.65,  288.65,
  288.6,     288.6,   288.6,   288.6,
  288.8,     288.8,   288.8,   288.8,
  288.95,    288.95,  288.95,  288.95,
  288.8,     288.8,   288.8,   288.8,
  288.75,    288.75,  288.75,  288.75,
  288.4,     288.4,   288.4,   288.4,
  287.7,     287.7,   287.7,   287.7,
  287.1,     287.1,   287.1,   287.1,
  286.7,     286.7,   286.7,   286.7,
  286.4,     286.4,   286.4,   286.4,
  286.15,    286.15,  286.15,  286.15,
  285.95,    285.95,  285.95,  285.95,
  285.7,     285.7,   285.7,   285.7,
  285.4,     285.4,   285.4,   285.4,
  285,       285,     285,     285,
  284.6,     284.6,   284.6,   284.6,
  284.35,    284.35,  284.35,  284.35,
  284.15,    284.15,  284.15,  284.15,
  283.85,    283.85,  283.85,  283.85,
  283.6,     283.6,   283.6,   283.6,
  283.55,    283.55,  283.55,  283.55,
  283.5,     283.5,   283.5,   283.5,
  283.4,     283.4,   283.4,   283.4,
  283.15,    283.15,  283.15,  283.15,
  282.8,     282.8,   282.8,   282.8,
  282.5,     282.5,   282.5,   282.5,
  282.2,     282.2,   282.2,   282.2,
  281.85,    281.85,  281.85,  281.85,
  281.55,    281.55,  281.55,  281.55,
  281.4,     281.4,   281.4,   281.4,
  281.25,    281.25,  281.25,  281.25,
  281.1,     281.1,   281.1,   281.1,
  281.1,     281.1,   281.1,   281.1,
  281.25,    281.25,  281.25,  281.25,
  281.6,     281.6,   281.6,   281.6,
  282.1,     282.1,   282.1,   282.1,
  282.8,     282.8,   282.8,   282.8,
  283.8,     283.8,   283.8,   283.8,
  285.05,    285.05,  285.05,  285.05,
  286.2,     286.2,   286.2,   286.2,
  287.2,     287.2,   287.2,   287.2,
  288.2,     288.2,   288.2,   288.2,
  288.95,    288.95,  288.95,  288.95,
  289.55,    289.55,  289.55,  289.55,
  290,       290,     290,     290,
  290.45,    290.45,  290.45,  290.45,
  290.9,     290.9,   290.9,   290.9,
  291.25,    291.25,  291.25,  291.25,
  291.55,    291.55,  291.55,  291.55,
  291.8,     291.8,   291.8,   291.8,
  292,       292,     292,     292,
  291.9,     291.9,   291.9,   291.9,
  291.5,     291.5,   291.5,   291.5,
  290.95,    290.95,  290.95,  290.95,
  290.15,    290.15,  290.15,  290.15,
  289.25,    289.25,  289.25,  289.25,
  288.5,     288.5,   288.5,   288.5,
  287.9,     287.9,   287.9,   287.9,
  287.4,     287.4,   287.4,   287.4,
  286.95,    286.95,  286.95,  286.95,
  286.45,    286.45,  286.45,  286.45,
  285.9,     285.9,   285.9,   285.9,
  285.6,     285.6,   285.6,   285.6,
  285.45,    285.45,  285.45,  285.45,
  285.2,     285.2,   285.2,   285.2,
  285,       285,     285,     285,
  284.9,     284.9,   284.9,   284.9,
  284.7,     284.7,   284.7,   284.7,
  284.4,     284.4,   284.4,   284.4,
  284.2,     284.2,   284.2,   284.2,
  284.05,    284.05,  284.05,  284.05,
  283.9,     283.9,   283.9,   283.9,
  283.95,    283.95,  283.95,  283.95,
  283.95,    283.95,  283.95,  283.95,
  283.65,    283.65,  283.65,  283.65,
  283.35,    283.35,  283.35,  283.35,
  283.15,    283.15,  283.15,  283.15,
  283,       283,     283,     283,
  282.9,     282.9,   282.9,   282.9,
  282.8,     282.8,   282.8,   282.8,
  282.7,     282.7,   282.7,   282.7,
  282.55,    282.55,  282.55,  282.55,
  282.45,    282.45,  282.45,  282.45,
  282.65,    282.65,  282.65,  282.65,
  283.25,    283.25,  283.25,  283.25,
  284.2,     284.2,   284.2,   284.2,
  285.15,    285.15,  285.15,  285.15,
  286,       286,     286,     286,
  286.9,     286.9,   286.9,   286.9,
  287.7,     287.7,   287.7,   287.7,
  288.55,    288.55,  288.55,  288.55,
  289.5,     289.5,   289.5,   289.5,
  290.2,     290.2,   290.2,   290.2,
  290.85,    290.85,  290.85,  290.85,
  291.6,     291.6,   291.6,   291.6,
  291.95,    291.95,  291.95,  291.95,
  291.95,    291.95,  291.95,  291.95,
  292,       292,     292,     292,
  292.1,     292.1,   292.1,   292.1,
  291.85,    291.85,  291.85,  291.85,
  291.35,    291.35,  291.35,  291.35,
  290.85,    290.85,  290.85,  290.85,
  290.45,    290.45,  290.45,  290.45,
  289.8,     289.8,   289.8,   289.8,
  289.05,    289.05,  289.05,  289.05,
  288.6,     288.6,   288.6,   288.6,
  288,       288,     288,     288,
  287.45,    287.45,  287.45,  287.45,
  287,       287,     287,     287,
  286.25,    286.25,  286.25,  286.25,
  285.55,    285.55,  285.55,  285.55,
  285.05,    285.05,  285.05,  285.05,
  284.5,     284.5,   284.5,   284.5,
  283.65,    283.65,  283.65,  283.65,
  282.75,    282.75,  282.75,  282.75,
  283,       283,     283,     283,
  283.95,    283.95,  283.95,  283.95,
  284.4,     284.4,   284.4,   284.4,
  284.75,    284.75,  284.75,  284.75,
  285.2,     285.2,   285.2,   285.2,
  285.4,     285.4,   285.4,   285.4,
  285.4,     285.4,   285.4,   285.4,
  285.3,     285.3,   285.3,   285.3,
  285.25,    285.25,  285.25,  285.25,
  285.2,     285.2,   285.2,   285.2,
  285.15,    285.15,  285.15,  285.15,
  285.15,    285.15,  285.15,  285.15,
  285.15,    285.15,  285.15,  285.15,
  285,       285,     285,     285,
  284.8,     284.8,   284.8,   284.8,
  284.7,     284.7,   284.7,   284.7,
  284.35,    284.35,  284.35,  284.35,
  283.85,    283.85,  283.85,  283.85,
  283.55,    283.55,  283.55,  283.55,
  283.35,    283.35,  283.35,  283.35,
  283.25,    283.25,  283.25,  283.25,
  283.3,     283.3,   283.3,   283.3,
  283.45,    283.45,  283.45,  283.45,
  283.6,     283.6,   283.6,   283.6,
  283.55,    283.55,  283.55,  283.55,
  283.45,    283.45,  283.45,  283.45,
  283.55,    283.55,  283.55,  283.55,
  283.55,    283.55,  283.55,  283.55,
  283.5,     283.5,   283.5,   283.5,
  283.55,    283.55,  283.55,  283.55,
  283.5,     283.5,   283.5,   283.5,
  283.15,    283.15,  283.15,  283.15,
  282.7,     282.7,   282.7,   282.7,
  282.3,     282.3,   282.3,   282.3,
  281.7,     281.7,   281.7,   281.7,
  280.85,    280.85,  280.85,  280.85,
  280.05,    280.05,  280.05,  280.05,
  279.4,     279.4,   279.4,   279.4,
  278.9,     278.9,   278.9,   278.9,
  278.5,     278.5,   278.5,   278.5,
  278.3,     278.3,   278.3,   278.3,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.2,     278.2,   278.2,   278.2,
  278,       278,     278,     278,
  277.95,    277.95,  277.95,  277.95,
  277.85,    277.85,  277.85,  277.85,
  277.6,     277.6,   277.6,   277.6,
  277.3,     277.3,   277.3,   277.3,
  277,       277,     277,     277,
  276.65,    276.65,  276.65,  276.65,
  276.25,    276.25,  276.25,  276.25,
  275.95,    275.95,  275.95,  275.95,
  275.75,    275.75,  275.75,  275.75,
  275.65,    275.65,  275.65,  275.65,
  275.7,     275.7,   275.7,   275.7,
  275.55,    275.55,  275.55,  275.55,
  275.2,     275.2,   275.2,   275.2,
  274.9,     274.9,   274.9,   274.9,
  274.6,     274.6,   274.6,   274.6,
  274.4,     274.4,   274.4,   274.4,
  274.35,    274.35,  274.35,  274.35,
  274.4,     274.4,   274.4,   274.4,
  274.5,     274.5,   274.5,   274.5,
  274.6,     274.6,   274.6,   274.6,
  274.85,    274.85,  274.85,  274.85,
  275.7,     275.7,   275.7,   275.7,
  277.05,    277.05,  277.05,  277.05,
  278.4,     278.4,   278.4,   278.4,
  279.4,     279.4,   279.4,   279.4,
  279.8,     279.8,   279.8,   279.8,
  280.2,     280.2,   280.2,   280.2,
  280.85,    280.85,  280.85,  280.85,
  281.3,     281.3,   281.3,   281.3,
  281.6,     281.6,   281.6,   281.6,
  281.85,    281.85,  281.85,  281.85,
  282,       282,     282,     282,
  282.15,    282.15,  282.15,  282.15,
  282.15,    282.15,  282.15,  282.15,
  282,       282,     282,     282,
  281.75,    281.75,  281.75,  281.75,
  281.35,    281.35,  281.35,  281.35,
  280.75,    280.75,  280.75,  280.75,
  280,       280,     280,     280,
  279.2,     279.2,   279.2,   279.2,
  278.45,    278.45,  278.45,  278.45,
  277.8,     277.8,   277.8,   277.8,
  277.1,     277.1,   277.1,   277.1,
  276.45,    276.45,  276.45,  276.45,
  276.2,     276.2,   276.2,   276.2,
  276.15,    276.15,  276.15,  276.15,
  275.95,    275.95,  275.95,  275.95,
  275.75,    275.75,  275.75,  275.75,
  275.8,     275.8,   275.8,   275.8,
  275.85,    275.85,  275.85,  275.85,
  275.6,     275.6,   275.6,   275.6,
  275.2,     275.2,   275.2,   275.2,
  274.7,     274.7,   274.7,   274.7,
  273.95,    273.95,  273.95,  273.95,
  273.45,    273.45,  273.45,  273.45,
  273.65,    273.65,  273.65,  273.65,
  273.5,     273.5,   273.5,   273.5,
  272.95,    272.95,  272.95,  272.95,
  272.7,     272.7,   272.7,   272.7,
  272.6,     272.6,   272.6,   272.6,
  272.6,     272.6,   272.6,   272.6,
  272.6,     272.6,   272.6,   272.6,
  272.65,    272.65,  272.65,  272.65,
  272.4,     272.4,   272.4,   272.4,
  272.15,    272.15,  272.15,  272.15,
  272.35,    272.35,  272.35,  272.35,
  272.4,     272.4,   272.4,   272.4,
  272.45,    272.45,  272.45,  272.45,
  273.4,     273.4,   273.4,   273.4,
  275.05,    275.05,  275.05,  275.05,
  276.35,    276.35,  276.35,  276.35,
  277.45,    277.45,  277.45,  277.45,
  278.65,    278.65,  278.65,  278.65,
  279.3,     279.3,   279.3,   279.3,
  279.85,    279.85,  279.85,  279.85,
  280.6,     280.6,   280.6,   280.6,
  281.2,     281.2,   281.2,   281.2,
  281.7,     281.7,   281.7,   281.7,
  282.1,     282.1,   282.1,   282.1,
  282.45,    282.45,  282.45,  282.45,
  282.8,     282.8,   282.8,   282.8,
  283.05,    283.05,  283.05,  283.05,
  283.15,    283.15,  283.15,  283.15,
  283,       283,     283,     283,
  282.45,    282.45,  282.45,  282.45,
  281.55,    281.55,  281.55,  281.55,
  280.25,    280.25,  280.25,  280.25,
  279.5,     279.5,   279.5,   279.5,
  279.45,    279.45,  279.45,  279.45,
  278.9,     278.9,   278.9,   278.9,
  277.6,     277.6,   277.6,   277.6,
  276.5,     276.5,   276.5,   276.5,
  276.15,    276.15,  276.15,  276.15,
  276.3,     276.3,   276.3,   276.3,
  276.05,    276.05,  276.05,  276.05,
  275.55,    275.55,  275.55,  275.55,
  275.15,    275.15,  275.15,  275.15,
  274.9,     274.9,   274.9,   274.9,
  274.85,    274.85,  274.85,  274.85,
  275,       275,     275,     275,
  275.45,    275.45,  275.45,  275.45,
  275.6,     275.6,   275.6,   275.6,
  275.8,     275.8,   275.8,   275.8,
  276,       276,     276,     276,
  275.95,    275.95,  275.95,  275.95,
  275.7,     275.7,   275.7,   275.7,
  275.7,     275.7,   275.7,   275.7,
  276.15,    276.15,  276.15,  276.15,
  276.3,     276.3,   276.3,   276.3,
  276.35,    276.35,  276.35,  276.35,
  276.35,    276.35,  276.35,  276.35,
  276.1,     276.1,   276.1,   276.1,
  276.2,     276.2,   276.2,   276.2,
  276.55,    276.55,  276.55,  276.55,
  276.75,    276.75,  276.75,  276.75,
  276.95,    276.95,  276.95,  276.95,
  277.1,     277.1,   277.1,   277.1,
  277.35,    277.35,  277.35,  277.35,
  277.9,     277.9,   277.9,   277.9,
  278.65,    278.65,  278.65,  278.65,
  279.65,    279.65,  279.65,  279.65,
  280.8,     280.8,   280.8,   280.8,
  281.9,     281.9,   281.9,   281.9,
  283.05,    283.05,  283.05,  283.05,
  283.5,     283.5,   283.5,   283.5,
  283.5,     283.5,   283.5,   283.5,
  283.45,    283.45,  283.45,  283.45,
  283.25,    283.25,  283.25,  283.25,
  283.3,     283.3,   283.3,   283.3,
  283.3,     283.3,   283.3,   283.3,
  283.4,     283.4,   283.4,   283.4,
  283.3,     283.3,   283.3,   283.3,
  282.85,    282.85,  282.85,  282.85,
  282.4,     282.4,   282.4,   282.4,
  281.85,    281.85,  281.85,  281.85,
  281.3,     281.3,   281.3,   281.3,
  280.95,    280.95,  280.95,  280.95,
  280.7,     280.7,   280.7,   280.7,
  280.35,    280.35,  280.35,  280.35,
  280.1,     280.1,   280.1,   280.1,
  280,       280,     280,     280,
  279.9,     279.9,   279.9,   279.9,
  279.8,     279.8,   279.8,   279.8,
  279.55,    279.55,  279.55,  279.55,
  279.35,    279.35,  279.35,  279.35,
  279.3,     279.3,   279.3,   279.3,
  279.15,    279.15,  279.15,  279.15,
  279.05,    279.05,  279.05,  279.05,
  279.2,     279.2,   279.2,   279.2,
  279.45,    279.45,  279.45,  279.45,
  279.5,     279.5,   279.5,   279.5,
  279.3,     279.3,   279.3,   279.3,
  278.85,    278.85,  278.85,  278.85,
  278.4,     278.4,   278.4,   278.4,
  277.95,    277.95,  277.95,  277.95,
  277.6,     277.6,   277.6,   277.6,
  277.65,    277.65,  277.65,  277.65,
  277.35,    277.35,  277.35,  277.35,
  276.8,     276.8,   276.8,   276.8,
  276.6,     276.6,   276.6,   276.6,
  276.35,    276.35,  276.35,  276.35,
  275.8,     275.8,   275.8,   275.8,
  275.6,     275.6,   275.6,   275.6,
  276,       276,     276,     276,
  276.75,    276.75,  276.75,  276.75,
  277.8,     277.8,   277.8,   277.8,
  278.6,     278.6,   278.6,   278.6,
  279.05,    279.05,  279.05,  279.05,
  279.6,     279.6,   279.6,   279.6,
  280.65,    280.65,  280.65,  280.65,
  281.4,     281.4,   281.4,   281.4,
  281.5,     281.5,   281.5,   281.5,
  281.7,     281.7,   281.7,   281.7,
  281.9,     281.9,   281.9,   281.9,
  282.1,     282.1,   282.1,   282.1,
  282.4,     282.4,   282.4,   282.4,
  282.35,    282.35,  282.35,  282.35,
  282,       282,     282,     282,
  281.85,    281.85,  281.85,  281.85,
  281.75,    281.75,  281.75,  281.75,
  281.45,    281.45,  281.45,  281.45,
  281,       281,     281,     281,
  280.5,     280.5,   280.5,   280.5,
  280,       280,     280,     280,
  279.5,     279.5,   279.5,   279.5,
  279.1,     279.1,   279.1,   279.1,
  278.85,    278.85,  278.85,  278.85,
  278.7,     278.7,   278.7,   278.7,
  278.5,     278.5,   278.5,   278.5,
  278.15,    278.15,  278.15,  278.15,
  277.85,    277.85,  277.85,  277.85,
  277.75,    277.75,  277.75,  277.75,
  277.75,    277.75,  277.75,  277.75,
  277.9,     277.9,   277.9,   277.9,
  278.1,     278.1,   278.1,   278.1,
  278.05,    278.05,  278.05,  278.05,
  277.8,     277.8,   277.8,   277.8,
  277.4,     277.4,   277.4,   277.4,
  276.95,    276.95,  276.95,  276.95,
  276.75,    276.75,  276.75,  276.75,
  276.65,    276.65,  276.65,  276.65,
  276.45,    276.45,  276.45,  276.45,
  276.25,    276.25,  276.25,  276.25,
  276.2,     276.2,   276.2,   276.2,
  276.25,    276.25,  276.25,  276.25,
  276.45,    276.45,  276.45,  276.45,
  276.9,     276.9,   276.9,   276.9,
  277.35,    277.35,  277.35,  277.35,
  277.75,    277.75,  277.75,  277.75,
  278.05,    278.05,  278.05,  278.05,
  278.25,    278.25,  278.25,  278.25,
  278.6,     278.6,   278.6,   278.6,
  279.15,    279.15,  279.15,  279.15,
  279.6,     279.6,   279.6,   279.6,
  280.1,     280.1,   280.1,   280.1,
  280.55,    280.55,  280.55,  280.55,
  281,       281,     281,     281,
  281.7,     281.7,   281.7,   281.7,
  282,       282,     282,     282,
  282.1,     282.1,   282.1,   282.1,
  282.55,    282.55,  282.55,  282.55,
  283.1,     283.1,   283.1,   283.1,
  283.35,    283.35,  283.35,  283.35,
  283.2,     283.2,   283.2,   283.2,
  283.05,    283.05,  283.05,  283.05,
  283.05,    283.05,  283.05,  283.05,
  283.1,     283.1,   283.1,   283.1,
  283.05,    283.05,  283.05,  283.05,
  282.6,     282.6,   282.6,   282.6,
  281.85,    281.85,  281.85,  281.85,
  281.3,     281.3,   281.3,   281.3,
  281.1,     281.1,   281.1,   281.1,
  281,       281,     281,     281,
  280.95,    280.95,  280.95,  280.95,
  280.9,     280.9,   280.9,   280.9,
  280.75,    280.75,  280.75,  280.75,
  280.5,     280.5,   280.5,   280.5,
  280.3,     280.3,   280.3,   280.3,
  280.25,    280.25,  280.25,  280.25,
  280.2,     280.2,   280.2,   280.2,
  280.15,    280.15,  280.15,  280.15,
  280.15,    280.15,  280.15,  280.15,
  280.15,    280.15,  280.15,  280.15,
  280.15,    280.15,  280.15,  280.15,
  279.9,     279.9,   279.9,   279.9,
  279.55,    279.55,  279.55,  279.55,
  279.35,    279.35,  279.35,  279.35,
  279.2,     279.2,   279.2,   279.2,
  279,       279,     279,     279,
  278.9,     278.9,   278.9,   278.9,
  278.75,    278.75,  278.75,  278.75,
  278.55,    278.55,  278.55,  278.55,
  278.55,    278.55,  278.55,  278.55,
  278.55,    278.55,  278.55,  278.55,
  278.6,     278.6,   278.6,   278.6,
  278.8,     278.8,   278.8,   278.8,
  279,       279,     279,     279,
  279.05,    279.05,  279.05,  279.05,
  279.05,    279.05,  279.05,  279.05,
  279.1,     279.1,   279.1,   279.1,
  279.35,    279.35,  279.35,  279.35,
  279.95,    279.95,  279.95,  279.95,
  280.65,    280.65,  280.65,  280.65,
  281.35,    281.35,  281.35,  281.35,
  282.05,    282.05,  282.05,  282.05,
  282.55,    282.55,  282.55,  282.55,
  283.05,    283.05,  283.05,  283.05,
  283.45,    283.45,  283.45,  283.45,
  283.65,    283.65,  283.65,  283.65,
  283.7,     283.7,   283.7,   283.7,
  283.7,     283.7,   283.7,   283.7,
  283.65,    283.65,  283.65,  283.65,
  283.15,    283.15,  283.15,  283.15,
  282.75,    282.75,  282.75,  282.75,
  282.5,     282.5,   282.5,   282.5,
  282.2,     282.2,   282.2,   282.2,
  282.05,    282.05,  282.05,  282.05,
  281.85,    281.85,  281.85,  281.85,
  281.65,    281.65,  281.65,  281.65,
  281.5,     281.5,   281.5,   281.5,
  281.3,     281.3,   281.3,   281.3,
  281.1,     281.1,   281.1,   281.1,
  281,       281,     281,     281,
  280.9,     280.9,   280.9,   280.9,
  280.8,     280.8,   280.8,   280.8,
  280.65,    280.65,  280.65,  280.65,
  280.45,    280.45,  280.45,  280.45,
  280.25,    280.25,  280.25,  280.25,
  280.05,    280.05,  280.05,  280.05,
  279.85,    279.85,  279.85,  279.85,
  279.65,    279.65,  279.65,  279.65,
  279.4,     279.4,   279.4,   279.4,
  279.05,    279.05,  279.05,  279.05,
  278.75,    278.75,  278.75,  278.75,
  278.55,    278.55,  278.55,  278.55,
  278.4,     278.4,   278.4,   278.4,
  278.3,     278.3,   278.3,   278.3,
  278.15,    278.15,  278.15,  278.15,
  277.95,    277.95,  277.95,  277.95,
  277.6,     277.6,   277.6,   277.6,
  277,       277,     277,     277,
  276.25,    276.25,  276.25,  276.25,
  275.55,    275.55,  275.55,  275.55,
  274.95,    274.95,  274.95,  274.95,
  274.5,     274.5,   274.5,   274.5,
  274.15,    274.15,  274.15,  274.15,
  273.8,     273.8,   273.8,   273.8,
  273.75,    273.75,  273.75,  273.75,
  274.05,    274.05,  274.05,  274.05,
  274.6,     274.6,   274.6,   274.6,
  275.25,    275.25,  275.25,  275.25,
  275.9,     275.9,   275.9,   275.9,
  276.6,     276.6,   276.6,   276.6,
  277.15,    277.15,  277.15,  277.15,
  277.5,     277.5,   277.5,   277.5,
  277.75,    277.75,  277.75,  277.75,
  277.95,    277.95,  277.95,  277.95,
  278.2,     278.2,   278.2,   278.2,
  278.4,     278.4,   278.4,   278.4,
  278.55,    278.55,  278.55,  278.55,
  278.65,    278.65,  278.65,  278.65,
  278.6,     278.6,   278.6,   278.6,
  278.55,    278.55,  278.55,  278.55,
  278.45,    278.45,  278.45,  278.45,
  278.1,     278.1,   278.1,   278.1,
  277.45,    277.45,  277.45,  277.45,
  276.6,     276.6,   276.6,   276.6,
  275.9,     275.9,   275.9,   275.9,
  275.55,    275.55,  275.55,  275.55,
  275.1,     275.1,   275.1,   275.1,
  274.55,    274.55,  274.55,  274.55,
  274.25,    274.25,  274.25,  274.25,
  274.05,    274.05,  274.05,  274.05,
  273.85,    273.85,  273.85,  273.85,
  273.65,    273.65,  273.65,  273.65,
  273.4,     273.4,   273.4,   273.4,
  273.1,     273.1,   273.1,   273.1,
  272.8,     272.8,   272.8,   272.8,
  272.45,    272.45,  272.45,  272.45,
  272.2,     272.2,   272.2,   272.2,
  272.05,    272.05,  272.05,  272.05,
  271.85,    271.85,  271.85,  271.85,
  271.6,     271.6,   271.6,   271.6,
  271.4,     271.4,   271.4,   271.4,
  271.4,     271.4,   271.4,   271.4,
  271.5,     271.5,   271.5,   271.5,
  271.5,     271.5,   271.5,   271.5,
  271.45,    271.45,  271.45,  271.45,
  271.35,    271.35,  271.35,  271.35,
  271.2,     271.2,   271.2,   271.2,
  271.15,    271.15,  271.15,  271.15,
  271.15,    271.15,  271.15,  271.15,
  271.1,     271.1,   271.1,   271.1,
  271.1,     271.1,   271.1,   271.1,
  271.05,    271.05,  271.05,  271.05,
  271.1,     271.1,   271.1,   271.1,
  271.75,    271.75,  271.75,  271.75,
  272.95,    272.95,  272.95,  272.95,
  274,       274,     274,     274,
  274.85,    274.85,  274.85,  274.85,
  275.9,     275.9,   275.9,   275.9,
  276.6,     276.6,   276.6,   276.6,
  276.95,    276.95,  276.95,  276.95,
  277.4,     277.4,   277.4,   277.4,
  277.8,     277.8,   277.8,   277.8,
  278.05,    278.05,  278.05,  278.05,
  278.35,    278.35,  278.35,  278.35,
  278.6,     278.6,   278.6,   278.6,
  278.75,    278.75,  278.75,  278.75,
  278.85,    278.85,  278.85,  278.85,
  278.85,    278.85,  278.85,  278.85,
  278.7,     278.7,   278.7,   278.7,
  278.2,     278.2,   278.2,   278.2,
  277.35,    277.35,  277.35,  277.35,
  276.35,    276.35,  276.35,  276.35,
  275.5,     275.5,   275.5,   275.5,
  275.1,     275.1,   275.1,   275.1,
  275.05,    275.05,  275.05,  275.05,
  274.8,     274.8,   274.8,   274.8,
  274.25,    274.25,  274.25,  274.25,
  273.6,     273.6,   273.6,   273.6,
  273.35,    273.35,  273.35,  273.35,
  273.4,     273.4,   273.4,   273.4,
  273.3,     273.3,   273.3,   273.3,
  272.95,    272.95,  272.95,  272.95,
  272.5,     272.5,   272.5,   272.5,
  272.15,    272.15,  272.15,  272.15,
  271.95,    271.95,  271.95,  271.95,
  272,       272,     272,     272,
  272.05,    272.05,  272.05,  272.05,
  271.75,    271.75,  271.75,  271.75,
  271.25,    271.25,  271.25,  271.25,
  270.95,    270.95,  270.95,  270.95,
  270.75,    270.75,  270.75,  270.75,
  270.4,     270.4,   270.4,   270.4,
  270.3,     270.3,   270.3,   270.3,
  270.3,     270.3,   270.3,   270.3,
  270.1,     270.1,   270.1,   270.1,
  270,       270,     270,     270,
  270,       270,     270,     270,
  270.05,    270.05,  270.05,  270.05,
  269.8,     269.8,   269.8,   269.8,
  269.85,    269.85,  269.85,  269.85,
  270.2,     270.2,   270.2,   270.2,
  270.7,     270.7,   270.7,   270.7,
  272,       272,     272,     272,
  273.4,     273.4,   273.4,   273.4,
  274.55,    274.55,  274.55,  274.55,
  275.95,    275.95,  275.95,  275.95,
  277.45,    277.45,  277.45,  277.45,
  278.4,     278.4,   278.4,   278.4,
  278.85,    278.85,  278.85,  278.85,
  279.3,     279.3,   279.3,   279.3,
  279.9,     279.9,   279.9,   279.9,
  280.35,    280.35,  280.35,  280.35,
  280.6,     280.6,   280.6,   280.6,
  280.85,    280.85,  280.85,  280.85,
  280.75,    280.75,  280.75,  280.75,
  280.5,     280.5,   280.5,   280.5,
  279.85,    279.85,  279.85,  279.85,
  278.7,     278.7,   278.7,   278.7,
  277.7,     277.7,   277.7,   277.7,
  276.9,     276.9,   276.9,   276.9,
  276.4,     276.4,   276.4,   276.4,
  276.15,    276.15,  276.15,  276.15,
  276.15,    276.15,  276.15,  276.15,
  276.1,     276.1,   276.1,   276.1,
  275.9,     275.9,   275.9,   275.9,
  275.7,     275.7,   275.7,   275.7,
  275.35,    275.35,  275.35,  275.35,
  274.55,    274.55,  274.55,  274.55,
  273.8,     273.8,   273.8,   273.8,
  273.7,     273.7,   273.7,   273.7,
  273.55,    273.55,  273.55,  273.55,
  273.4,     273.4,   273.4,   273.4,
  273.8,     273.8,   273.8,   273.8,
  274.25,    274.25,  274.25,  274.25,
  274.2,     274.2,   274.2,   274.2,
  274,       274,     274,     274,
  273.8,     273.8,   273.8,   273.8,
  273.5,     273.5,   273.5,   273.5,
  273.45,    273.45,  273.45,  273.45,
  273.6,     273.6,   273.6,   273.6,
  273.8,     273.8,   273.8,   273.8,
  274.05,    274.05,  274.05,  274.05,
  273.75,    273.75,  273.75,  273.75,
  273.4,     273.4,   273.4,   273.4,
  273.25,    273.25,  273.25,  273.25,
  273.25,    273.25,  273.25,  273.25,
  273.45,    273.45,  273.45,  273.45,
  273.65,    273.65,  273.65,  273.65,
  273.9,     273.9,   273.9,   273.9,
  274.05,    274.05,  274.05,  274.05,
  274.5,     274.5,   274.5,   274.5,
  275.25,    275.25,  275.25,  275.25,
  276.05,    276.05,  276.05,  276.05,
  277.1,     277.1,   277.1,   277.1,
  278.4,     278.4,   278.4,   278.4,
  279.75,    279.75,  279.75,  279.75,
  281.1,     281.1,   281.1,   281.1,
  282.35,    282.35,  282.35,  282.35,
  283.1,     283.1,   283.1,   283.1,
  283.35,    283.35,  283.35,  283.35,
  283.7,     283.7,   283.7,   283.7,
  283.85,    283.85,  283.85,  283.85,
  283.55,    283.55,  283.55,  283.55,
  283.15,    283.15,  283.15,  283.15,
  282.7,     282.7,   282.7,   282.7,
  282.1,     282.1,   282.1,   282.1,
  281.15,    281.15,  281.15,  281.15,
  280.05,    280.05,  280.05,  280.05,
  279.15,    279.15,  279.15,  279.15,
  278.25,    278.25,  278.25,  278.25,
  277.75,    277.75,  277.75,  277.75,
  277.65,    277.65,  277.65,  277.65,
  277.55,    277.55,  277.55,  277.55,
  277.6,     277.6,   277.6,   277.6,
  277.95,    277.95,  277.95,  277.95,
  278.35,    278.35,  278.35,  278.35,
  278.2,     278.2,   278.2,   278.2,
  277.85,    277.85,  277.85,  277.85,
  277.65,    277.65,  277.65,  277.65,
  277.45,    277.45,  277.45,  277.45,
  277.4,     277.4,   277.4,   277.4,
  277.25,    277.25,  277.25,  277.25,
  276.95,    276.95,  276.95,  276.95,
  276.55,    276.55,  276.55,  276.55,
  275.9,     275.9,   275.9,   275.9,
  275.65,    275.65,  275.65,  275.65,
  275.7,     275.7,   275.7,   275.7,
  275.55,    275.55,  275.55,  275.55,
  275.25,    275.25,  275.25,  275.25,
  274.25,    274.25,  274.25,  274.25,
  273.3,     273.3,   273.3,   273.3,
  273.2,     273.2,   273.2,   273.2,
  273.85,    273.85,  273.85,  273.85,
  274.7,     274.7,   274.7,   274.7,
  274.9,     274.9,   274.9,   274.9,
  275.25,    275.25,  275.25,  275.25,
  276,       276,     276,     276,
  276.7,     276.7,   276.7,   276.7,
  277.5,     277.5,   277.5,   277.5,
  278.35,    278.35,  278.35,  278.35,
  279.1,     279.1,   279.1,   279.1,
  279.9,     279.9,   279.9,   279.9,
  280.65,    280.65,  280.65,  280.65,
  281.3,     281.3,   281.3,   281.3,
  282,       282,     282,     282,
  282.7,     282.7,   282.7,   282.7,
  283.35,    283.35,  283.35,  283.35,
  283.8,     283.8,   283.8,   283.8,
  284,       284,     284,     284,
  284.05,    284.05,  284.05,  284.05,
  284,       284,     284,     284,
  283.8,     283.8,   283.8,   283.8,
  283.45,    283.45,  283.45,  283.45,
  282.95,    282.95,  282.95,  282.95,
  282.2,     282.2,   282.2,   282.2,
  281.25,    281.25,  281.25,  281.25,
  280.5,     280.5,   280.5,   280.5,
  280.1,     280.1,   280.1,   280.1,
  279.55,    279.55,  279.55,  279.55,
  279,       279,     279,     279,
  278.85,    278.85,  278.85,  278.85,
  278.6,     278.6,   278.6,   278.6,
  278.1,     278.1,   278.1,   278.1,
  277.2,     277.2,   277.2,   277.2,
  276.35,    276.35,  276.35,  276.35,
  276.1,     276.1,   276.1,   276.1,
  275.85,    275.85,  275.85,  275.85,
  275.4,     275.4,   275.4,   275.4,
  275.1,     275.1,   275.1,   275.1,
  275.05,    275.05,  275.05,  275.05,
  274.95,    274.95,  274.95,  274.95,
  274.75,    274.75,  274.75,  274.75,
  274.6,     274.6,   274.6,   274.6,
  274.6,     274.6,   274.6,   274.6,
  274.7,     274.7,   274.7,   274.7,
  274.75,    274.75,  274.75,  274.75,
  274.75,    274.75,  274.75,  274.75,
  274.75,    274.75,  274.75,  274.75,
  274.75,    274.75,  274.75,  274.75,
  274.8,     274.8,   274.8,   274.8,
  274.95,    274.95,  274.95,  274.95,
  275.1,     275.1,   275.1,   275.1,
  275.25,    275.25,  275.25,  275.25,
  275.35,    275.35,  275.35,  275.35,
  275.3,     275.3,   275.3,   275.3,
  275.25,    275.25,  275.25,  275.25,
  275.3,     275.3,   275.3,   275.3,
  275.4,     275.4,   275.4,   275.4,
  275.5,     275.5,   275.5,   275.5,
  275.65,    275.65,  275.65,  275.65,
  275.85,    275.85,  275.85,  275.85,
  276,       276,     276,     276,
  276.05,    276.05,  276.05,  276.05,
  276.1,     276.1,   276.1,   276.1,
  276.15,    276.15,  276.15,  276.15,
  276.35,    276.35,  276.35,  276.35,
  276.55,    276.55,  276.55,  276.55,
  276.75,    276.75,  276.75,  276.75,
  277.05,    277.05,  277.05,  277.05,
  277,       277,     277,     277,
  276.8,     276.8,   276.8,   276.8,
  276.55,    276.55,  276.55,  276.55,
  275.85,    275.85,  275.85,  275.85,
  274.95,    274.95,  274.95,  274.95,
  274.35,    274.35,  274.35,  274.35,
  273.8,     273.8,   273.8,   273.8,
  273.15,    273.15,  273.15,  273.15,
  272.75,    272.75,  272.75,  272.75,
  272.5,     272.5,   272.5,   272.5,
  272.1,     272.1,   272.1,   272.1,
  271.7,     271.7,   271.7,   271.7,
  271.55,    271.55,  271.55,  271.55,
  271.4,     271.4,   271.4,   271.4,
  271,       271,     271,     271,
  270.45,    270.45,  270.45,  270.45,
  270,       270,     270,     270,
  269.75,    269.75,  269.75,  269.75,
  269.7,     269.7,   269.7,   269.7,
  269.9,     269.9,   269.9,   269.9,
  270.2,     270.2,   270.2,   270.2,
  270.5,     270.5,   270.5,   270.5,
  270.75,    270.75,  270.75,  270.75,
  271.2,     271.2,   271.2,   271.2,
  271.65,    271.65,  271.65,  271.65,
  271.8,     271.8,   271.8,   271.8,
  271.9,     271.9,   271.9,   271.9,
  271.95,    271.95,  271.95,  271.95,
  271.95,    271.95,  271.95,  271.95,
  272,       272,     272,     272,
  272.05,    272.05,  272.05,  272.05,
  272,       272,     272,     272,
  271.9,     271.9,   271.9,   271.9,
  271.85,    271.85,  271.85,  271.85,
  271.9,     271.9,   271.9,   271.9,
  271.8,     271.8,   271.8,   271.8,
  271.7,     271.7,   271.7,   271.7,
  271.95,    271.95,  271.95,  271.95,
  272.3,     272.3,   272.3,   272.3,
  272.65,    272.65,  272.65,  272.65,
  273.25,    273.25,  273.25,  273.25,
  273.95,    273.95,  273.95,  273.95,
  274.55,    274.55,  274.55,  274.55,
  275,       275,     275,     275,
  275.25,    275.25,  275.25,  275.25,
  275.4,     275.4,   275.4,   275.4,
  275.6,     275.6,   275.6,   275.6,
  275.85,    275.85,  275.85,  275.85,
  276,       276,     276,     276,
  276.15,    276.15,  276.15,  276.15,
  276.35,    276.35,  276.35,  276.35,
  276.5,     276.5,   276.5,   276.5,
  276.6,     276.6,   276.6,   276.6,
  276.65,    276.65,  276.65,  276.65,
  276.55,    276.55,  276.55,  276.55,
  276.4,     276.4,   276.4,   276.4,
  276.35,    276.35,  276.35,  276.35,
  276.35,    276.35,  276.35,  276.35,
  276.35,    276.35,  276.35,  276.35,
  276.4,     276.4,   276.4,   276.4,
  276.45,    276.45,  276.45,  276.45,
  276.45,    276.45,  276.45,  276.45,
  276.45,    276.45,  276.45,  276.45,
  276.5,     276.5,   276.5,   276.5,
  276.5,     276.5,   276.5,   276.5,
  276.5,     276.5,   276.5,   276.5,
  276.55,    276.55,  276.55,  276.55,
  276.6,     276.6,   276.6,   276.6,
  276.65,    276.65,  276.65,  276.65,
  276.6,     276.6,   276.6,   276.6,
  276.55,    276.55,  276.55,  276.55,
  276.6,     276.6,   276.6,   276.6,
  276.65,    276.65,  276.65,  276.65,
  276.65,    276.65,  276.65,  276.65,
  276.65,    276.65,  276.65,  276.65,
  276.65,    276.65,  276.65,  276.65,
  276.65,    276.65,  276.65,  276.65,
  276.65,    276.65,  276.65,  276.65,
  276.65,    276.65,  276.65,  276.65,
  276.65,    276.65,  276.65,  276.65,
  276.65,    276.65,  276.65,  276.65,
  276.7,     276.7,   276.7,   276.7,
  276.8,     276.8,   276.8,   276.8,
  277.05,    277.05,  277.05,  277.05,
  277.5,     277.5,   277.5,   277.5,
  278.1,     278.1,   278.1,   278.1,
  278.7,     278.7,   278.7,   278.7,
  279.35,    279.35,  279.35,  279.35,
  280.4,     280.4,   280.4,   280.4,
  281.3,     281.3,   281.3,   281.3,
  281.35,    281.35,  281.35,  281.35,
  281.1,     281.1,   281.1,   281.1,
  280.85,    280.85,  280.85,  280.85,
  280.5,     280.5,   280.5,   280.5,
  280.25,    280.25,  280.25,  280.25,
  280.2,     280.2,   280.2,   280.2,
  280.3,     280.3,   280.3,   280.3,
  280.35,    280.35,  280.35,  280.35,
  280.3,     280.3,   280.3,   280.3,
  280.15,    280.15,  280.15,  280.15,
  280,       280,     280,     280,
  279.8,     279.8,   279.8,   279.8,
  279.55,    279.55,  279.55,  279.55,
  279.2,     279.2,   279.2,   279.2,
  278.75,    278.75,  278.75,  278.75,
  278.3,     278.3,   278.3,   278.3,
  277.95,    277.95,  277.95,  277.95,
  277.7,     277.7,   277.7,   277.7,
  277.35,    277.35,  277.35,  277.35,
  276.9,     276.9,   276.9,   276.9,
  276.5,     276.5,   276.5,   276.5,
  276.2,     276.2,   276.2,   276.2,
  275.9,     275.9,   275.9,   275.9,
  275.6,     275.6,   275.6,   275.6,
  275.35,    275.35,  275.35,  275.35,
  275.15,    275.15,  275.15,  275.15,
  274.95,    274.95,  274.95,  274.95,
  274.75,    274.75,  274.75,  274.75,
  274.55,    274.55,  274.55,  274.55,
  274.4,     274.4,   274.4,   274.4,
  274.25,    274.25,  274.25,  274.25,
  274.05,    274.05,  274.05,  274.05,
  273.9,     273.9,   273.9,   273.9,
  273.8,     273.8,   273.8,   273.8,
  273.7,     273.7,   273.7,   273.7,
  273.55,    273.55,  273.55,  273.55,
  273.35,    273.35,  273.35,  273.35,
  273.1,     273.1,   273.1,   273.1,
  272.95,    272.95,  272.95,  272.95,
  273,       273,     273,     273,
  273.25,    273.25,  273.25,  273.25,
  273.75,    273.75,  273.75,  273.75,
  274.55,    274.55,  274.55,  274.55,
  275.65,    275.65,  275.65,  275.65,
  276.7,     276.7,   276.7,   276.7,
  277.55,    277.55,  277.55,  277.55,
  278.2,     278.2,   278.2,   278.2,
  278.85,    278.85,  278.85,  278.85,
  279.4,     279.4,   279.4,   279.4,
  279.8,     279.8,   279.8,   279.8,
  280.25,    280.25,  280.25,  280.25,
  280.55,    280.55,  280.55,  280.55,
  280.7,     280.7,   280.7,   280.7,
  280.75,    280.75,  280.75,  280.75,
  280.65,    280.65,  280.65,  280.65,
  280.4,     280.4,   280.4,   280.4,
  279.95,    279.95,  279.95,  279.95,
  279.35,    279.35,  279.35,  279.35,
  278.9,     278.9,   278.9,   278.9,
  278.75,    278.75,  278.75,  278.75,
  278.65,    278.65,  278.65,  278.65,
  278.5,     278.5,   278.5,   278.5,
  278.25,    278.25,  278.25,  278.25,
  278.05,    278.05,  278.05,  278.05,
  278.05,    278.05,  278.05,  278.05,
  278.15,    278.15,  278.15,  278.15,
  278.4,     278.4,   278.4,   278.4,
  278.75,    278.75,  278.75,  278.75,
  279.05,    279.05,  279.05,  279.05,
  279.15,    279.15,  279.15,  279.15,
  279.05,    279.05,  279.05,  279.05,
  278.7,     278.7,   278.7,   278.7,
  278.2,     278.2,   278.2,   278.2,
  277.95,    277.95,  277.95,  277.95,
  278.05,    278.05,  278.05,  278.05,
  278.2,     278.2,   278.2,   278.2,
  278.35,    278.35,  278.35,  278.35,
  278.6,     278.6,   278.6,   278.6,
  278.85,    278.85,  278.85,  278.85,
  279.1,     279.1,   279.1,   279.1,
  279.35,    279.35,  279.35,  279.35,
  279.55,    279.55,  279.55,  279.55,
  279.85,    279.85,  279.85,  279.85,
  280.2,     280.2,   280.2,   280.2,
  280.5,     280.5,   280.5,   280.5,
  280.85,    280.85,  280.85,  280.85,
  281.1,     281.1,   281.1,   281.1,
  281.35,    281.35,  281.35,  281.35,
  281.7,     281.7,   281.7,   281.7,
  282.05,    282.05,  282.05,  282.05,
  282.6,     282.6,   282.6,   282.6,
  283.2,     283.2,   283.2,   283.2,
  283.55,    283.55,  283.55,  283.55,
  283.95,    283.95,  283.95,  283.95,
  284.6,     284.6,   284.6,   284.6,
  285.35,    285.35,  285.35,  285.35,
  286.2,     286.2,   286.2,   286.2,
  286.8,     286.8,   286.8,   286.8,
  286.95,    286.95,  286.95,  286.95,
  287,       287,     287,     287,
  287.2,     287.2,   287.2,   287.2,
  287.2,     287.2,   287.2,   287.2,
  287,       287,     287,     287,
  286.85,    286.85,  286.85,  286.85,
  286.55,    286.55,  286.55,  286.55,
  285.95,    285.95,  285.95,  285.95,
  285.2,     285.2,   285.2,   285.2,
  284.55,    284.55,  284.55,  284.55,
  284.15,    284.15,  284.15,  284.15,
  283.9,     283.9,   283.9,   283.9,
  283.65,    283.65,  283.65,  283.65,
  283.4,     283.4,   283.4,   283.4,
  283.05,    283.05,  283.05,  283.05,
  282.75,    282.75,  282.75,  282.75,
  282.6,     282.6,   282.6,   282.6,
  282.5,     282.5,   282.5,   282.5,
  282.45,    282.45,  282.45,  282.45,
  282.6,     282.6,   282.6,   282.6,
  282.85,    282.85,  282.85,  282.85,
  283,       283,     283,     283,
  283.1,     283.1,   283.1,   283.1,
  283.1,     283.1,   283.1,   283.1,
  283.05,    283.05,  283.05,  283.05,
  283.1,     283.1,   283.1,   283.1,
  283.2,     283.2,   283.2,   283.2,
  283.35,    283.35,  283.35,  283.35,
  283.35,    283.35,  283.35,  283.35,
  283.25,    283.25,  283.25,  283.25,
  283.35,    283.35,  283.35,  283.35,
  283.5,     283.5,   283.5,   283.5,
  283.55,    283.55,  283.55,  283.55,
  283.5,     283.5,   283.5,   283.5,
  283.4,     283.4,   283.4,   283.4,
  283.25,    283.25,  283.25,  283.25,
  283.15,    283.15,  283.15,  283.15,
  283.2,     283.2,   283.2,   283.2,
  283.25,    283.25,  283.25,  283.25,
  283.35,    283.35,  283.35,  283.35,
  283.55,    283.55,  283.55,  283.55,
  283.85,    283.85,  283.85,  283.85,
  284.3,     284.3,   284.3,   284.3,
  284.65,    284.65,  284.65,  284.65,
  284.9,     284.9,   284.9,   284.9,
  285.15,    285.15,  285.15,  285.15,
  285.35,    285.35,  285.35,  285.35,
  285.45,    285.45,  285.45,  285.45,
  285.6,     285.6,   285.6,   285.6,
  285.85,    285.85,  285.85,  285.85,
  285.95,    285.95,  285.95,  285.95,
  285.9,     285.9,   285.9,   285.9,
  285.9,     285.9,   285.9,   285.9,
  285.9,     285.9,   285.9,   285.9,
  285.5,     285.5,   285.5,   285.5,
  284.85,    284.85,  284.85,  284.85,
  284.4,     284.4,   284.4,   284.4,
  284,       284,     284,     284,
  283.5,     283.5,   283.5,   283.5,
  283.15,    283.15,  283.15,  283.15,
  282.95,    282.95,  282.95,  282.95,
  282.9,     282.9,   282.9,   282.9,
  282.95,    282.95,  282.95,  282.95,
  283,       283,     283,     283,
  283.1,     283.1,   283.1,   283.1,
  283.1,     283.1,   283.1,   283.1,
  283.05,    283.05,  283.05,  283.05,
  283.3,     283.3,   283.3,   283.3,
  283.65,    283.65,  283.65,  283.65,
  283.8,     283.8,   283.8,   283.8,
  283.75,    283.75,  283.75,  283.75,
  283.6,     283.6,   283.6,   283.6,
  283.5,     283.5,   283.5,   283.5,
  283.45,    283.45,  283.45,  283.45,
  283.55,    283.55,  283.55,  283.55,
  283.65,    283.65,  283.65,  283.65,
  283.65,    283.65,  283.65,  283.65,
  283.8,     283.8,   283.8,   283.8,
  284.25,    284.25,  284.25,  284.25,
  284.9,     284.9,   284.9,   284.9,
  285.45,    285.45,  285.45,  285.45,
  285.7,     285.7,   285.7,   285.7,
  285.6,     285.6,   285.6,   285.6,
  284.65,    284.65,  284.65,  284.65,
  283.6,     283.6,   283.6,   283.6,
  283.4,     283.4,   283.4,   283.4,
  283.5,     283.5,   283.5,   283.5,
  283.55,    283.55,  283.55,  283.55,
  283.5,     283.5,   283.5,   283.5,
  283.25,    283.25,  283.25,  283.25,
  283.15,    283.15,  283.15,  283.15,
  283.35,    283.35,  283.35,  283.35,
  283.25,    283.25,  283.25,  283.25,
  283,       283,     283,     283,
  282.95,    282.95,  282.95,  282.95,
  282.9,     282.9,   282.9,   282.9,
  282.9,     282.9,   282.9,   282.9,
  283,       283,     283,     283,
  283.05,    283.05,  283.05,  283.05,
  283.05,    283.05,  283.05,  283.05,
  283.05,    283.05,  283.05,  283.05,
  283.1,     283.1,   283.1,   283.1,
  283.2,     283.2,   283.2,   283.2,
  283.3,     283.3,   283.3,   283.3,
  283.35,    283.35,  283.35,  283.35,
  283.4,     283.4,   283.4,   283.4,
  283.5,     283.5,   283.5,   283.5,
  283.6,     283.6,   283.6,   283.6,
  283.6,     283.6,   283.6,   283.6,
  283.6,     283.6,   283.6,   283.6,
  283.5,     283.5,   283.5,   283.5,
  283.1,     283.1,   283.1,   283.1,
  282.65,    282.65,  282.65,  282.65,
  282.45,    282.45,  282.45,  282.45,
  282.4,     282.4,   282.4,   282.4,
  282.2,     282.2,   282.2,   282.2,
  281.7,     281.7,   281.7,   281.7,
  281.1,     281.1,   281.1,   281.1,
  280.85,    280.85,  280.85,  280.85,
  281.05,    281.05,  281.05,  281.05,
  281.6,     281.6,   281.6,   281.6,
  282.1,     282.1,   282.1,   282.1,
  282,       282,     282,     282,
  281.7,     281.7,   281.7,   281.7,
  281.75,    281.75,  281.75,  281.75,
  281.75,    281.75,  281.75,  281.75,
  281.7,     281.7,   281.7,   281.7,
  281.8,     281.8,   281.8,   281.8,
  281.9,     281.9,   281.9,   281.9,
  282.05,    282.05,  282.05,  282.05,
  282.15,    282.15,  282.15,  282.15,
  282.05,    282.05,  282.05,  282.05,
  281.85,    281.85,  281.85,  281.85,
  282.05,    282.05,  282.05,  282.05,
  282.5,     282.5,   282.5,   282.5,
  282.85,    282.85,  282.85,  282.85,
  283,       283,     283,     283,
  282.9,     282.9,   282.9,   282.9,
  282.9,     282.9,   282.9,   282.9,
  283.05,    283.05,  283.05,  283.05,
  283.35,    283.35,  283.35,  283.35,
  283.65,    283.65,  283.65,  283.65,
  284,       284,     284,     284,
  284.4,     284.4,   284.4,   284.4,
  284.6,     284.6,   284.6,   284.6,
  284.7,     284.7,   284.7,   284.7,
  284.95,    284.95,  284.95,  284.95,
  285.2,     285.2,   285.2,   285.2,
  285.15,    285.15,  285.15,  285.15,
  284.9,     284.9,   284.9,   284.9,
  284.55,    284.55,  284.55,  284.55,
  284.2,     284.2,   284.2,   284.2,
  283.95,    283.95,  283.95,  283.95,
  283.85,    283.85,  283.85,  283.85,
  283.8,     283.8,   283.8,   283.8,
  283.6,     283.6,   283.6,   283.6,
  283.25,    283.25,  283.25,  283.25,
  282.8,     282.8,   282.8,   282.8,
  282.5,     282.5,   282.5,   282.5,
  282.4,     282.4,   282.4,   282.4,
  282.3,     282.3,   282.3,   282.3,
  282.25,    282.25,  282.25,  282.25,
  282.3,     282.3,   282.3,   282.3,
  282.65,    282.65,  282.65,  282.65,
  283.15,    283.15,  283.15,  283.15,
  283.25,    283.25,  283.25,  283.25,
  283.15,    283.15,  283.15,  283.15,
  283.3,     283.3,   283.3,   283.3,
  282.95,    282.95,  282.95,  282.95,
  282.2,     282.2,   282.2,   282.2,
  281.9,     281.9,   281.9,   281.9,
  281.85,    281.85,  281.85,  281.85,
  281.95,    281.95,  281.95,  281.95,
  282.1,     282.1,   282.1,   282.1,
  282.2,     282.2,   282.2,   282.2,
  282.3,     282.3,   282.3,   282.3,
  282.45,    282.45,  282.45,  282.45,
  282.55,    282.55,  282.55,  282.55,
  282.5,     282.5,   282.5,   282.5,
  282.3,     282.3,   282.3,   282.3,
  281.6,     281.6,   281.6,   281.6,
  281,       281,     281,     281,
  280.9,     280.9,   280.9,   280.9,
  281.1,     281.1,   281.1,   281.1,
  281.75,    281.75,  281.75,  281.75,
  282.4,     282.4,   282.4,   282.4,
  282.85,    282.85,  282.85,  282.85,
  283.2,     283.2,   283.2,   283.2,
  283.6,     283.6,   283.6,   283.6,
  284.05,    284.05,  284.05,  284.05,
  284.25,    284.25,  284.25,  284.25,
  284.35,    284.35,  284.35,  284.35,
  284.45,    284.45,  284.45,  284.45,
  284.45,    284.45,  284.45,  284.45,
  284.55,    284.55,  284.55,  284.55,
  284.75,    284.75,  284.75,  284.75,
  284.7,     284.7,   284.7,   284.7,
  284.15,    284.15,  284.15,  284.15,
  283.55,    283.55,  283.55,  283.55,
  283.2,     283.2,   283.2,   283.2,
  282.9,     282.9,   282.9,   282.9,
  282.65,    282.65,  282.65,  282.65,
  282.55,    282.55,  282.55,  282.55,
  282.55,    282.55,  282.55,  282.55,
  282.4,     282.4,   282.4,   282.4,
  282.1,     282.1,   282.1,   282.1,
  281.9,     281.9,   281.9,   281.9,
  281.75,    281.75,  281.75,  281.75,
  281.5,     281.5,   281.5,   281.5,
  281.25,    281.25,  281.25,  281.25,
  281,       281,     281,     281,
  280.85,    280.85,  280.85,  280.85,
  281.3,     281.3,   281.3,   281.3,
  281.7,     281.7,   281.7,   281.7,
  281.65,    281.65,  281.65,  281.65,
  281.55,    281.55,  281.55,  281.55,
  281.35,    281.35,  281.35,  281.35,
  281.4,     281.4,   281.4,   281.4,
  281.45,    281.45,  281.45,  281.45,
  281.15,    281.15,  281.15,  281.15,
  280.95,    280.95,  280.95,  280.95,
  280.85,    280.85,  280.85,  280.85,
  280.7,     280.7,   280.7,   280.7,
  280.55,    280.55,  280.55,  280.55,
  280.35,    280.35,  280.35,  280.35,
  280.2,     280.2,   280.2,   280.2,
  280.25,    280.25,  280.25,  280.25,
  280.65,    280.65,  280.65,  280.65,
  281,       281,     281,     281,
  281.05,    281.05,  281.05,  281.05,
  281.2,     281.2,   281.2,   281.2,
  281.55,    281.55,  281.55,  281.55,
  281.9,     281.9,   281.9,   281.9,
  282.15,    282.15,  282.15,  282.15,
  282.4,     282.4,   282.4,   282.4,
  282.7,     282.7,   282.7,   282.7,
  283.15,    283.15,  283.15,  283.15,
  283.4,     283.4,   283.4,   283.4,
  283.55,    283.55,  283.55,  283.55,
  283.8,     283.8,   283.8,   283.8,
  284.05,    284.05,  284.05,  284.05,
  284.5,     284.5,   284.5,   284.5,
  284.65,    284.65,  284.65,  284.65,
  284.35,    284.35,  284.35,  284.35,
  284.1,     284.1,   284.1,   284.1,
  284,       284,     284,     284,
  283.85,    283.85,  283.85,  283.85,
  283.55,    283.55,  283.55,  283.55,
  282.95,    282.95,  282.95,  282.95,
  281.95,    281.95,  281.95,  281.95,
  281.3,     281.3,   281.3,   281.3,
  281.2,     281.2,   281.2,   281.2,
  281.15,    281.15,  281.15,  281.15,
  281.2,     281.2,   281.2,   281.2,
  281.3,     281.3,   281.3,   281.3,
  281.3,     281.3,   281.3,   281.3,
  281.15,    281.15,  281.15,  281.15,
  281,       281,     281,     281,
  280.95,    280.95,  280.95,  280.95,
  280.85,    280.85,  280.85,  280.85,
  280.6,     280.6,   280.6,   280.6,
  280.65,    280.65,  280.65,  280.65,
  280.85,    280.85,  280.85,  280.85,
  280.8,     280.8,   280.8,   280.8,
  280.85,    280.85,  280.85,  280.85,
  281,       281,     281,     281,
  281,       281,     281,     281,
  281,       281,     281,     281,
  281,       281,     281,     281,
  280.9,     280.9,   280.9,   280.9,
  280.75,    280.75,  280.75,  280.75,
  280.6,     280.6,   280.6,   280.6,
  280.35,    280.35,  280.35,  280.35,
  279.85,    279.85,  279.85,  279.85,
  279.4,     279.4,   279.4,   279.4,
  279.2,     279.2,   279.2,   279.2,
  279.05,    279.05,  279.05,  279.05,
  278.85,    278.85,  278.85,  278.85,
  279,       279,     279,     279,
  279.55,    279.55,  279.55,  279.55,
  280.15,    280.15,  280.15,  280.15,
  280.7,     280.7,   280.7,   280.7,
  281.15,    281.15,  281.15,  281.15,
  281.35,    281.35,  281.35,  281.35,
  281.4,     281.4,   281.4,   281.4,
  281.6,     281.6,   281.6,   281.6,
  281.65,    281.65,  281.65,  281.65,
  281.25,    281.25,  281.25,  281.25,
  280.65,    280.65,  280.65,  280.65,
  280.15,    280.15,  280.15,  280.15,
  279.65,    279.65,  279.65,  279.65,
  279.25,    279.25,  279.25,  279.25,
  279.1,     279.1,   279.1,   279.1,
  279.05,    279.05,  279.05,  279.05,
  279.05,    279.05,  279.05,  279.05,
  279.1,     279.1,   279.1,   279.1,
  279.2,     279.2,   279.2,   279.2,
  279.35,    279.35,  279.35,  279.35,
  279.55,    279.55,  279.55,  279.55,
  279.6,     279.6,   279.6,   279.6,
  279.55,    279.55,  279.55,  279.55,
  279.55,    279.55,  279.55,  279.55,
  279.4,     279.4,   279.4,   279.4,
  279.2,     279.2,   279.2,   279.2,
  279.3,     279.3,   279.3,   279.3,
  279.6,     279.6,   279.6,   279.6,
  279.9,     279.9,   279.9,   279.9,
  280.05,    280.05,  280.05,  280.05,
  279.9,     279.9,   279.9,   279.9,
  279.5,     279.5,   279.5,   279.5,
  279.1,     279.1,   279.1,   279.1,
  278.75,    278.75,  278.75,  278.75,
  278.35,    278.35,  278.35,  278.35,
  278.05,    278.05,  278.05,  278.05,
  277.95,    277.95,  277.95,  277.95,
  278.1,     278.1,   278.1,   278.1,
  278,       278,     278,     278,
  277.65,    277.65,  277.65,  277.65,
  277.55,    277.55,  277.55,  277.55,
  277.45,    277.45,  277.45,  277.45,
  277.35,    277.35,  277.35,  277.35,
  277,       277,     277,     277,
  276.6,     276.6,   276.6,   276.6,
  276.75,    276.75,  276.75,  276.75,
  277.35,    277.35,  277.35,  277.35,
  277,       277,     277,     277,
  276.4,     276.4,   276.4,   276.4,
  276,       276,     276,     276,
  275.8,     275.8,   275.8,   275.8,
  276.7,     276.7,   276.7,   276.7,
  277.5,     277.5,   277.5,   277.5,
  278.25,    278.25,  278.25,  278.25,
  279.25,    279.25,  279.25,  279.25,
  279.95,    279.95,  279.95,  279.95,
  280.35,    280.35,  280.35,  280.35,
  280.75,    280.75,  280.75,  280.75,
  281.05,    281.05,  281.05,  281.05,
  281.2,     281.2,   281.2,   281.2,
  281.3,     281.3,   281.3,   281.3,
  281.3,     281.3,   281.3,   281.3,
  281.1,     281.1,   281.1,   281.1,
  280.75,    280.75,  280.75,  280.75,
  280.35,    280.35,  280.35,  280.35,
  280,       280,     280,     280,
  279.7,     279.7,   279.7,   279.7,
  279.5,     279.5,   279.5,   279.5,
  279.3,     279.3,   279.3,   279.3,
  278.9,     278.9,   278.9,   278.9,
  278.3,     278.3,   278.3,   278.3,
  277.7,     277.7,   277.7,   277.7,
  277.35,    277.35,  277.35,  277.35,
  277.3,     277.3,   277.3,   277.3,
  277.45,    277.45,  277.45,  277.45,
  277.55,    277.55,  277.55,  277.55,
  277.65,    277.65,  277.65,  277.65,
  277.7,     277.7,   277.7,   277.7,
  277.55,    277.55,  277.55,  277.55,
  277.5,     277.5,   277.5,   277.5,
  277.65,    277.65,  277.65,  277.65,
  277.8,     277.8,   277.8,   277.8,
  277.85,    277.85,  277.85,  277.85,
  277.85,    277.85,  277.85,  277.85,
  277.9,     277.9,   277.9,   277.9,
  278.05,    278.05,  278.05,  278.05,
  278.05,    278.05,  278.05,  278.05,
  277.8,     277.8,   277.8,   277.8,
  277.6,     277.6,   277.6,   277.6,
  277.45,    277.45,  277.45,  277.45,
  277.3,     277.3,   277.3,   277.3,
  277.2,     277.2,   277.2,   277.2,
  277.2,     277.2,   277.2,   277.2,
  277.2,     277.2,   277.2,   277.2,
  277.15,    277.15,  277.15,  277.15,
  277.2,     277.2,   277.2,   277.2,
  277.15,    277.15,  277.15,  277.15,
  277.1,     277.1,   277.1,   277.1,
  277.3,     277.3,   277.3,   277.3,
  277.55,    277.55,  277.55,  277.55,
  277.65,    277.65,  277.65,  277.65,
  277.6,     277.6,   277.6,   277.6,
  277.65,    277.65,  277.65,  277.65,
  277.85,    277.85,  277.85,  277.85,
  278.05,    278.05,  278.05,  278.05,
  278.25,    278.25,  278.25,  278.25,
  278.45,    278.45,  278.45,  278.45,
  278.5,     278.5,   278.5,   278.5,
  278.45,    278.45,  278.45,  278.45,
  278.4,     278.4,   278.4,   278.4,
  278.4,     278.4,   278.4,   278.4,
  278.5,     278.5,   278.5,   278.5,
  278.6,     278.6,   278.6,   278.6,
  278.6,     278.6,   278.6,   278.6,
  278.5,     278.5,   278.5,   278.5,
  278.35,    278.35,  278.35,  278.35,
  278.2,     278.2,   278.2,   278.2,
  278.25,    278.25,  278.25,  278.25,
  278.45,    278.45,  278.45,  278.45,
  278.65,    278.65,  278.65,  278.65,
  278.8,     278.8,   278.8,   278.8,
  278.8,     278.8,   278.8,   278.8,
  278.75,    278.75,  278.75,  278.75,
  278.6,     278.6,   278.6,   278.6,
  278.4,     278.4,   278.4,   278.4,
  278.35,    278.35,  278.35,  278.35,
  278.3,     278.3,   278.3,   278.3,
  278.3,     278.3,   278.3,   278.3,
  278.2,     278.2,   278.2,   278.2,
  277.95,    277.95,  277.95,  277.95,
  277.6,     277.6,   277.6,   277.6,
  277.1,     277.1,   277.1,   277.1,
  276.95,    276.95,  276.95,  276.95,
  277.2,     277.2,   277.2,   277.2,
  277.35,    277.35,  277.35,  277.35,
  277.3,     277.3,   277.3,   277.3,
  277.3,     277.3,   277.3,   277.3,
  277.3,     277.3,   277.3,   277.3,
  277.1,     277.1,   277.1,   277.1,
  276.9,     276.9,   276.9,   276.9,
  276.75,    276.75,  276.75,  276.75,
  276.55,    276.55,  276.55,  276.55,
  276.45,    276.45,  276.45,  276.45,
  276.45,    276.45,  276.45,  276.45,
  276.5,     276.5,   276.5,   276.5,
  276.7,     276.7,   276.7,   276.7,
  277.15,    277.15,  277.15,  277.15,
  277.75,    277.75,  277.75,  277.75,
  278.6,     278.6,   278.6,   278.6,
  279.4,     279.4,   279.4,   279.4,
  279.75,    279.75,  279.75,  279.75,
  279.95,    279.95,  279.95,  279.95,
  280,       280,     280,     280,
  279.9,     279.9,   279.9,   279.9,
  279.95,    279.95,  279.95,  279.95,
  280.15,    280.15,  280.15,  280.15,
  280.3,     280.3,   280.3,   280.3,
  280.3,     280.3,   280.3,   280.3,
  280.3,     280.3,   280.3,   280.3,
  280.4,     280.4,   280.4,   280.4,
  280.4,     280.4,   280.4,   280.4,
  280.35,    280.35,  280.35,  280.35,
  280.35,    280.35,  280.35,  280.35,
  280.35,    280.35,  280.35,  280.35,
  280.3,     280.3,   280.3,   280.3,
  280.25,    280.25,  280.25,  280.25,
  280,       280,     280,     280,
  279.75,    279.75,  279.75,  279.75,
  279.7,     279.7,   279.7,   279.7,
  279.45,    279.45,  279.45,  279.45,
  279.25,    279.25,  279.25,  279.25,
  279.45,    279.45,  279.45,  279.45,
  279.85,    279.85,  279.85,  279.85,
  280.1,     280.1,   280.1,   280.1,
  280.2,     280.2,   280.2,   280.2,
  280.25,    280.25,  280.25,  280.25,
  280.25,    280.25,  280.25,  280.25,
  280.35,    280.35,  280.35,  280.35,
  280.55,    280.55,  280.55,  280.55,
  280.6,     280.6,   280.6,   280.6,
  280.6,     280.6,   280.6,   280.6,
  280.55,    280.55,  280.55,  280.55,
  280.35,    280.35,  280.35,  280.35,
  280.2,     280.2,   280.2,   280.2,
  280.05,    280.05,  280.05,  280.05,
  279.95,    279.95,  279.95,  279.95,
  279.95,    279.95,  279.95,  279.95,
  279.95,    279.95,  279.95,  279.95,
  280.05,    280.05,  280.05,  280.05,
  280.2,     280.2,   280.2,   280.2,
  280.3,     280.3,   280.3,   280.3,
  280.45,    280.45,  280.45,  280.45,
  280.6,     280.6,   280.6,   280.6,
  280.7,     280.7,   280.7,   280.7,
  280.8,     280.8,   280.8,   280.8,
  280.9,     280.9,   280.9,   280.9,
  281.05,    281.05,  281.05,  281.05,
  281.2,     281.2,   281.2,   281.2,
  281.35,    281.35,  281.35,  281.35,
  281.5,     281.5,   281.5,   281.5,
  281.6,     281.6,   281.6,   281.6,
  281.75,    281.75,  281.75,  281.75,
  281.9,     281.9,   281.9,   281.9,
  282.05,    282.05,  282.05,  282.05,
  282.25,    282.25,  282.25,  282.25,
  282.4,     282.4,   282.4,   282.4,
  282.5,     282.5,   282.5,   282.5,
  282.55,    282.55,  282.55,  282.55,
  282.6,     282.6,   282.6,   282.6,
  282.65,    282.65,  282.65,  282.65,
  282.7,     282.7,   282.7,   282.7,
  282.8,     282.8,   282.8,   282.8,
  282.9,     282.9,   282.9,   282.9,
  282.95,    282.95,  282.95,  282.95,
  282.95,    282.95,  282.95,  282.95,
  283,       283,     283,     283,
  283.05,    283.05,  283.05,  283.05,
  283.05,    283.05,  283.05,  283.05,
  283.1,     283.1,   283.1,   283.1,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  283.2,     283.2,   283.2,   283.2,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.3,     283.3,   283.3,   283.3,
  283.35,    283.35,  283.35,  283.35,
  283.35,    283.35,  283.35,  283.35,
  283.3,     283.3,   283.3,   283.3,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.3,     283.3,   283.3,   283.3,
  283.3,     283.3,   283.3,   283.3,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.2,     283.2,   283.2,   283.2,
  283.2,     283.2,   283.2,   283.2,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.25,    283.25,  283.25,  283.25,
  283.3,     283.3,   283.3,   283.3,
  283.45,    283.45,  283.45,  283.45,
  283.55,    283.55,  283.55,  283.55,
  283.55,    283.55,  283.55,  283.55,
  283.5,     283.5,   283.5,   283.5,
  283.45,    283.45,  283.45,  283.45,
  283.4,     283.4,   283.4,   283.4,
  283.35,    283.35,  283.35,  283.35,
  283.4,     283.4,   283.4,   283.4,
  283.45,    283.45,  283.45,  283.45,
  283.5,     283.5,   283.5,   283.5,
  283.5,     283.5,   283.5,   283.5,
  283.35,    283.35,  283.35,  283.35,
  283.2,     283.2,   283.2,   283.2,
  283.05,    283.05,  283.05,  283.05,
  282.9,     282.9,   282.9,   282.9,
  282.65,    282.65,  282.65,  282.65,
  282.3,     282.3,   282.3,   282.3,
  281.95,    281.95,  281.95,  281.95,
  281.65,    281.65,  281.65,  281.65,
  281.45,    281.45,  281.45,  281.45,
  281.4,     281.4,   281.4,   281.4,
  281.3,     281.3,   281.3,   281.3,
  281.05,    281.05,  281.05,  281.05,
  280.9,     280.9,   280.9,   280.9,
  280.7,     280.7,   280.7,   280.7,
  280.35,    280.35,  280.35,  280.35,
  279.85,    279.85,  279.85,  279.85,
  279.35,    279.35,  279.35,  279.35,
  278.95,    278.95,  278.95,  278.95,
  278.6,     278.6,   278.6,   278.6,
  278.35,    278.35,  278.35,  278.35,
  278.3,     278.3,   278.3,   278.3,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.3,     278.3,   278.3,   278.3,
  278.2,     278.2,   278.2,   278.2,
  278.1,     278.1,   278.1,   278.1,
  277.95,    277.95,  277.95,  277.95,
  277.7,     277.7,   277.7,   277.7,
  277.45,    277.45,  277.45,  277.45,
  277.25,    277.25,  277.25,  277.25,
  277.15,    277.15,  277.15,  277.15,
  277.15,    277.15,  277.15,  277.15,
  277.15,    277.15,  277.15,  277.15,
  277.3,     277.3,   277.3,   277.3,
  277.7,     277.7,   277.7,   277.7,
  278.25,    278.25,  278.25,  278.25,
  278.8,     278.8,   278.8,   278.8,
  279.2,     279.2,   279.2,   279.2,
  279.55,    279.55,  279.55,  279.55,
  280,       280,     280,     280,
  280.6,     280.6,   280.6,   280.6,
  281.1,     281.1,   281.1,   281.1,
  281.35,    281.35,  281.35,  281.35,
  281.4,     281.4,   281.4,   281.4,
  281.2,     281.2,   281.2,   281.2,
  281,       281,     281,     281,
  280.75,    280.75,  280.75,  280.75,
  280.2,     280.2,   280.2,   280.2,
  279.7,     279.7,   279.7,   279.7,
  279.3,     279.3,   279.3,   279.3,
  278.95,    278.95,  278.95,  278.95,
  278.8,     278.8,   278.8,   278.8,
  278.65,    278.65,  278.65,  278.65,
  278.35,    278.35,  278.35,  278.35,
  278,       278,     278,     278,
  277.65,    277.65,  277.65,  277.65,
  277.4,     277.4,   277.4,   277.4,
  277.35,    277.35,  277.35,  277.35,
  277.1,     277.1,   277.1,   277.1,
  276.8,     276.8,   276.8,   276.8,
  276.65,    276.65,  276.65,  276.65,
  276.4,     276.4,   276.4,   276.4,
  276.1,     276.1,   276.1,   276.1,
  275.7,     275.7,   275.7,   275.7,
  275.3,     275.3,   275.3,   275.3,
  275,       275,     275,     275,
  274.7,     274.7,   274.7,   274.7,
  274.5,     274.5,   274.5,   274.5,
  274.45,    274.45,  274.45,  274.45,
  274.45,    274.45,  274.45,  274.45,
  274.5,     274.5,   274.5,   274.5,
  274.6,     274.6,   274.6,   274.6,
  274.75,    274.75,  274.75,  274.75,
  274.9,     274.9,   274.9,   274.9,
  274.9,     274.9,   274.9,   274.9,
  274.85,    274.85,  274.85,  274.85,
  274.9,     274.9,   274.9,   274.9,
  274.9,     274.9,   274.9,   274.9,
  274.8,     274.8,   274.8,   274.8,
  274.9,     274.9,   274.9,   274.9,
  275.25,    275.25,  275.25,  275.25,
  275.8,     275.8,   275.8,   275.8,
  276.55,    276.55,  276.55,  276.55,
  277.4,     277.4,   277.4,   277.4,
  278.15,    278.15,  278.15,  278.15,
  278.65,    278.65,  278.65,  278.65,
  279,       279,     279,     279,
  279.3,     279.3,   279.3,   279.3,
  279.7,     279.7,   279.7,   279.7,
  280.15,    280.15,  280.15,  280.15,
  280.55,    280.55,  280.55,  280.55,
  280.85,    280.85,  280.85,  280.85,
  281,       281,     281,     281,
  281.05,    281.05,  281.05,  281.05,
  280.9,     280.9,   280.9,   280.9,
  280.5,     280.5,   280.5,   280.5,
  279.9,     279.9,   279.9,   279.9,
  279.4,     279.4,   279.4,   279.4,
  279.1,     279.1,   279.1,   279.1,
  278.8,     278.8,   278.8,   278.8,
  278.4,     278.4,   278.4,   278.4,
  277.85,    277.85,  277.85,  277.85,
  277.4,     277.4,   277.4,   277.4,
  277.15,    277.15,  277.15,  277.15,
  276.95,    276.95,  276.95,  276.95,
  276.75,    276.75,  276.75,  276.75,
  276.6,     276.6,   276.6,   276.6,
  276.45,    276.45,  276.45,  276.45,
  276.3,     276.3,   276.3,   276.3,
  276.15,    276.15,  276.15,  276.15,
  275.9,     275.9,   275.9,   275.9,
  275.7,     275.7,   275.7,   275.7,
  275.55,    275.55,  275.55,  275.55,
  275.35,    275.35,  275.35,  275.35,
  275.35,    275.35,  275.35,  275.35,
  275.6,     275.6,   275.6,   275.6,
  275.85,    275.85,  275.85,  275.85,
  275.95,    275.95,  275.95,  275.95,
  276.05,    276.05,  276.05,  276.05,
  276,       276,     276,     276,
  275.65,    275.65,  275.65,  275.65,
  275.1,     275.1,   275.1,   275.1,
  274.45,    274.45,  274.45,  274.45,
  273.95,    273.95,  273.95,  273.95,
  273.6,     273.6,   273.6,   273.6,
  273.4,     273.4,   273.4,   273.4,
  273.4,     273.4,   273.4,   273.4,
  273.6,     273.6,   273.6,   273.6,
  273.7,     273.7,   273.7,   273.7,
  273.7,     273.7,   273.7,   273.7,
  274.05,    274.05,  274.05,  274.05,
  274.65,    274.65,  274.65,  274.65,
  275.15,    275.15,  275.15,  275.15,
  275.6,     275.6,   275.6,   275.6,
  276.2,     276.2,   276.2,   276.2,
  276.85,    276.85,  276.85,  276.85,
  277.35,    277.35,  277.35,  277.35,
  277.75,    277.75,  277.75,  277.75,
  278.1,     278.1,   278.1,   278.1,
  278.2,     278.2,   278.2,   278.2,
  278.15,    278.15,  278.15,  278.15,
  278.1,     278.1,   278.1,   278.1,
  277.9,     277.9,   277.9,   277.9,
  277.4,     277.4,   277.4,   277.4,
  276.75,    276.75,  276.75,  276.75,
  276.15,    276.15,  276.15,  276.15,
  275.6,     275.6,   275.6,   275.6,
  275.2,     275.2,   275.2,   275.2,
  275,       275,     275,     275,
  274.8,     274.8,   274.8,   274.8,
  274.5,     274.5,   274.5,   274.5,
  274.4,     274.4,   274.4,   274.4,
  274.45,    274.45,  274.45,  274.45,
  274.35,    274.35,  274.35,  274.35,
  274,       274,     274,     274,
  273.3,     273.3,   273.3,   273.3,
  272.7,     272.7,   272.7,   272.7,
  272.6,     272.6,   272.6,   272.6,
  272.8,     272.8,   272.8,   272.8,
  273.05,    273.05,  273.05,  273.05,
  273.15,    273.15,  273.15,  273.15,
  272.95,    272.95,  272.95,  272.95,
  272.6,     272.6,   272.6,   272.6,
  272.45,    272.45,  272.45,  272.45,
  272.45,    272.45,  272.45,  272.45,
  272.6,     272.6,   272.6,   272.6,
  272.8,     272.8,   272.8,   272.8,
  272.85,    272.85,  272.85,  272.85,
  272.85,    272.85,  272.85,  272.85,
  272.85,    272.85,  272.85,  272.85,
  272.9,     272.9,   272.9,   272.9,
  273,       273,     273,     273,
  273.05,    273.05,  273.05,  273.05,
  273.05,    273.05,  273.05,  273.05,
  272.8,     272.8,   272.8,   272.8,
  272.45,    272.45,  272.45,  272.45,
  272.4,     272.4,   272.4,   272.4,
  272.5,     272.5,   272.5,   272.5,
  272.8,     272.8,   272.8,   272.8,
  273.2,     273.2,   273.2,   273.2,
  273.15,    273.15,  273.15,  273.15,
  273.05,    273.05,  273.05,  273.05,
  273.35,    273.35,  273.35,  273.35,
  273.75,    273.75,  273.75,  273.75,
  274.3,     274.3,   274.3,   274.3,
  275.1,     275.1,   275.1,   275.1,
  275.75,    275.75,  275.75,  275.75,
  275.95,    275.95,  275.95,  275.95,
  276,       276,     276,     276,
  276.2,     276.2,   276.2,   276.2,
  276.4,     276.4,   276.4,   276.4,
  276.45,    276.45,  276.45,  276.45,
  276.5,     276.5,   276.5,   276.5,
  276.7,     276.7,   276.7,   276.7,
  277.1,     277.1,   277.1,   277.1,
  277.45,    277.45,  277.45,  277.45,
  277.5,     277.5,   277.5,   277.5,
  277.35,    277.35,  277.35,  277.35,
  277.4,     277.4,   277.4,   277.4,
  277.65,    277.65,  277.65,  277.65,
  277.8,     277.8,   277.8,   277.8,
  277.85,    277.85,  277.85,  277.85,
  277.95,    277.95,  277.95,  277.95,
  278.15,    278.15,  278.15,  278.15,
  278.25,    278.25,  278.25,  278.25,
  278.3,     278.3,   278.3,   278.3,
  278.4,     278.4,   278.4,   278.4,
  278.55,    278.55,  278.55,  278.55,
  278.7,     278.7,   278.7,   278.7,
  278.6,     278.6,   278.6,   278.6,
  278.5,     278.5,   278.5,   278.5,
  278.55,    278.55,  278.55,  278.55,
  278.6,     278.6,   278.6,   278.6,
  278.95,    278.95,  278.95,  278.95,
  279.5,     279.5,   279.5,   279.5,
  279.9,     279.9,   279.9,   279.9,
  280.1,     280.1,   280.1,   280.1,
  280.25,    280.25,  280.25,  280.25,
  280.4,     280.4,   280.4,   280.4,
  280.35,    280.35,  280.35,  280.35,
  280.15,    280.15,  280.15,  280.15,
  280,       280,     280,     280,
  280,       280,     280,     280,
  280.15,    280.15,  280.15,  280.15,
  280.3,     280.3,   280.3,   280.3,
  280.45,    280.45,  280.45,  280.45,
  280.7,     280.7,   280.7,   280.7,
  280.95,    280.95,  280.95,  280.95,
  281.2,     281.2,   281.2,   281.2,
  281.5,     281.5,   281.5,   281.5,
  281.8,     281.8,   281.8,   281.8,
  282,       282,     282,     282,
  282.05,    282.05,  282.05,  282.05,
  282.1,     282.1,   282.1,   282.1,
  282.1,     282.1,   282.1,   282.1,
  282,       282,     282,     282,
  281.9,     281.9,   281.9,   281.9,
  281.8,     281.8,   281.8,   281.8,
  281.7,     281.7,   281.7,   281.7,
  281.65,    281.65,  281.65,  281.65,
  281.55,    281.55,  281.55,  281.55,
  281.35,    281.35,  281.35,  281.35,
  281.25,    281.25,  281.25,  281.25,
  281.2,     281.2,   281.2,   281.2,
  281,       281,     281,     281,
  280.8,     280.8,   280.8,   280.8,
  280.75,    280.75,  280.75,  280.75,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.5,     280.5,   280.5,   280.5,
  280.3,     280.3,   280.3,   280.3,
  280.25,    280.25,  280.25,  280.25,
  280.25,    280.25,  280.25,  280.25,
  280.2,     280.2,   280.2,   280.2,
  280.2,     280.2,   280.2,   280.2,
  280.25,    280.25,  280.25,  280.25,
  280.25,    280.25,  280.25,  280.25,
  280.35,    280.35,  280.35,  280.35,
  280.6,     280.6,   280.6,   280.6,
  280.55,    280.55,  280.55,  280.55,
  280.3,     280.3,   280.3,   280.3,
  280.2,     280.2,   280.2,   280.2,
  280.05,    280.05,  280.05,  280.05,
  280.15,    280.15,  280.15,  280.15,
  280.2,     280.2,   280.2,   280.2,
  279.9,     279.9,   279.9,   279.9,
  279.65,    279.65,  279.65,  279.65,
  279.5,     279.5,   279.5,   279.5,
  279.45,    279.45,  279.45,  279.45,
  279.45,    279.45,  279.45,  279.45,
  279.45,    279.45,  279.45,  279.45,
  279.4,     279.4,   279.4,   279.4,
  279.3,     279.3,   279.3,   279.3,
  279.25,    279.25,  279.25,  279.25,
  279.3,     279.3,   279.3,   279.3,
  279.4,     279.4,   279.4,   279.4,
  279.75,    279.75,  279.75,  279.75,
  280.2,     280.2,   280.2,   280.2,
  280.5,     280.5,   280.5,   280.5,
  280.75,    280.75,  280.75,  280.75,
  280.85,    280.85,  280.85,  280.85,
  280.85,    280.85,  280.85,  280.85,
  280.85,    280.85,  280.85,  280.85,
  280.9,     280.9,   280.9,   280.9,
  280.85,    280.85,  280.85,  280.85,
  280.65,    280.65,  280.65,  280.65,
  280.4,     280.4,   280.4,   280.4,
  280.05,    280.05,  280.05,  280.05,
  279.55,    279.55,  279.55,  279.55,
  279.05,    279.05,  279.05,  279.05,
  278.65,    278.65,  278.65,  278.65,
  278.45,    278.45,  278.45,  278.45,
  278.55,    278.55,  278.55,  278.55,
  278.55,    278.55,  278.55,  278.55,
  278.4,     278.4,   278.4,   278.4,
  278.4,     278.4,   278.4,   278.4,
  278.45,    278.45,  278.45,  278.45,
  278.5,     278.5,   278.5,   278.5,
  278.5,     278.5,   278.5,   278.5,
  278.45,    278.45,  278.45,  278.45,
  278.45,    278.45,  278.45,  278.45,
  278.4,     278.4,   278.4,   278.4,
  278.4,     278.4,   278.4,   278.4,
  278.35,    278.35,  278.35,  278.35,
  278.1,     278.1,   278.1,   278.1,
  277.9,     277.9,   277.9,   277.9,
  277.75,    277.75,  277.75,  277.75,
  277.65,    277.65,  277.65,  277.65,
  277.65,    277.65,  277.65,  277.65,
  277.65,    277.65,  277.65,  277.65,
  277.6,     277.6,   277.6,   277.6,
  277.45,    277.45,  277.45,  277.45,
  277.35,    277.35,  277.35,  277.35,
  277.35,    277.35,  277.35,  277.35,
  277.35,    277.35,  277.35,  277.35,
  277.4,     277.4,   277.4,   277.4,
  277.5,     277.5,   277.5,   277.5,
  277.6,     277.6,   277.6,   277.6,
  277.65,    277.65,  277.65,  277.65,
  277.65,    277.65,  277.65,  277.65,
  277.7,     277.7,   277.7,   277.7,
  277.75,    277.75,  277.75,  277.75,
  277.8,     277.8,   277.8,   277.8,
  277.9,     277.9,   277.9,   277.9,
  278.05,    278.05,  278.05,  278.05,
  278.25,    278.25,  278.25,  278.25,
  278.5,     278.5,   278.5,   278.5,
  278.7,     278.7,   278.7,   278.7,
  278.8,     278.8,   278.8,   278.8,
  278.95,    278.95,  278.95,  278.95,
  279.1,     279.1,   279.1,   279.1,
  279.15,    279.15,  279.15,  279.15,
  279.15,    279.15,  279.15,  279.15,
  279.15,    279.15,  279.15,  279.15,
  279.15,    279.15,  279.15,  279.15,
  279.15,    279.15,  279.15,  279.15,
  279.1,     279.1,   279.1,   279.1,
  279,       279,     279,     279,
  278.9,     278.9,   278.9,   278.9,
  278.75,    278.75,  278.75,  278.75,
  278.55,    278.55,  278.55,  278.55,
  278.4,     278.4,   278.4,   278.4,
  278.3,     278.3,   278.3,   278.3,
  278.25,    278.25,  278.25,  278.25,
  278.25,    278.25,  278.25,  278.25,
  278.2,     278.2,   278.2,   278.2,
  278.05,    278.05,  278.05,  278.05,
  277.95,    277.95,  277.95,  277.95,
  277.95,    277.95,  277.95,  277.95,
  277.9,     277.9,   277.9,   277.9,
  277.75,    277.75,  277.75,  277.75,
  277.6,     277.6,   277.6,   277.6,
  277.55,    277.55,  277.55,  277.55,
  277.5,     277.5,   277.5,   277.5,
  277.45,    277.45,  277.45,  277.45,
  277.45,    277.45,  277.45,  277.45,
  277.3,     277.3,   277.3,   277.3,
  277.05,    277.05,  277.05,  277.05,
  276.8,     276.8,   276.8,   276.8,
  276.4,     276.4,   276.4,   276.4,
  275.8,     275.8,   275.8,   275.8,
  275.2,     275.2,   275.2,   275.2,
  274.9,     274.9,   274.9,   274.9,
  274.9,     274.9,   274.9,   274.9,
  274.95,    274.95,  274.95,  274.95,
  274.9,     274.9,   274.9,   274.9,
  274.8,     274.8,   274.8,   274.8,
  274.65,    274.65,  274.65,  274.65,
  274.45,    274.45,  274.45,  274.45,
  274.4,     274.4,   274.4,   274.4,
  274.55,    274.55,  274.55,  274.55,
  274.85,    274.85,  274.85,  274.85,
  275.25,    275.25,  275.25,  275.25,
  275.5,     275.5,   275.5,   275.5,
  275.55,    275.55,  275.55,  275.55,
  275.6,     275.6,   275.6,   275.6,
  275.7,     275.7,   275.7,   275.7,
  275.8,     275.8,   275.8,   275.8,
  275.85,    275.85,  275.85,  275.85,
  275.75,    275.75,  275.75,  275.75,
  275.65,    275.65,  275.65,  275.65,
  275.55,    275.55,  275.55,  275.55,
  275.4,     275.4,   275.4,   275.4,
  275.35,    275.35,  275.35,  275.35,
  275.15,    275.15,  275.15,  275.15,
  274.85,    274.85,  274.85,  274.85,
  274.75,    274.75,  274.75,  274.75,
  274.85,    274.85,  274.85,  274.85,
  274.9,     274.9,   274.9,   274.9,
  274.75,    274.75,  274.75,  274.75,
  274.7,     274.7,   274.7,   274.7,
  274.7,     274.7,   274.7,   274.7,
  274.55,    274.55,  274.55,  274.55,
  274.45,    274.45,  274.45,  274.45,
  274.45,    274.45,  274.45,  274.45,
  274.5,     274.5,   274.5,   274.5,
  274.55,    274.55,  274.55,  274.55,
  274.5,     274.5,   274.5,   274.5,
  274.4,     274.4,   274.4,   274.4,
  274.25,    274.25,  274.25,  274.25,
  274.1,     274.1,   274.1,   274.1,
  274,       274,     274,     274,
  273.85,    273.85,  273.85,  273.85,
  273.7,     273.7,   273.7,   273.7,
  273.6,     273.6,   273.6,   273.6,
  273.5,     273.5,   273.5,   273.5,
  273.45,    273.45,  273.45,  273.45,
  273.4,     273.4,   273.4,   273.4,
  273.35,    273.35,  273.35,  273.35,
  273.4,     273.4,   273.4,   273.4,
  273.5,     273.5,   273.5,   273.5,
  273.6,     273.6,   273.6,   273.6,
  273.7,     273.7,   273.7,   273.7,
  273.75,    273.75,  273.75,  273.75,
  273.85,    273.85,  273.85,  273.85,
  274.1,     274.1,   274.1,   274.1,
  274.35,    274.35,  274.35,  274.35,
  274.45,    274.45,  274.45,  274.45,
  274.45,    274.45,  274.45,  274.45,
  274.7,     274.7,   274.7,   274.7,
  275.4,     275.4,   275.4,   275.4,
  276.15,    276.15,  276.15,  276.15,
  276.55,    276.55,  276.55,  276.55,
  276.8,     276.8,   276.8,   276.8,
  277.1,     277.1,   277.1,   277.1,
  277.4,     277.4,   277.4,   277.4,
  277.85,    277.85,  277.85,  277.85,
  278.25,    278.25,  278.25,  278.25,
  278.35,    278.35,  278.35,  278.35,
  278.3,     278.3,   278.3,   278.3,
  278.05,    278.05,  278.05,  278.05,
  277.7,     277.7,   277.7,   277.7,
  277.45,    277.45,  277.45,  277.45,
  277.15,    277.15,  277.15,  277.15,
  276.8,     276.8,   276.8,   276.8,
  276.55,    276.55,  276.55,  276.55,
  276.5,     276.5,   276.5,   276.5,
  276.4,     276.4,   276.4,   276.4,
  276.2,     276.2,   276.2,   276.2,
  276.05,    276.05,  276.05,  276.05,
  276.1,     276.1,   276.1,   276.1,
  276.35,    276.35,  276.35,  276.35,
  276.3,     276.3,   276.3,   276.3,
  276.2,     276.2,   276.2,   276.2,
  276.35,    276.35,  276.35,  276.35,
  276.05,    276.05,  276.05,  276.05,
  275.35,    275.35,  275.35,  275.35,
  274.95,    274.95,  274.95,  274.95,
  274.85,    274.85,  274.85,  274.85,
  274.75,    274.75,  274.75,  274.75,
  274.5,     274.5,   274.5,   274.5,
  274.25,    274.25,  274.25,  274.25,
  274,       274,     274,     274,
  273.85,    273.85,  273.85,  273.85,
  274,       274,     274,     274,
  274.25,    274.25,  274.25,  274.25,
  274.3,     274.3,   274.3,   274.3,
  274.2,     274.2,   274.2,   274.2,
  274.05,    274.05,  274.05,  274.05,
  273.85,    273.85,  273.85,  273.85,
  273.75,    273.75,  273.75,  273.75,
  273.8,     273.8,   273.8,   273.8,
  273.75,    273.75,  273.75,  273.75,
  273.65,    273.65,  273.65,  273.65,
  273.6,     273.6,   273.6,   273.6,
  273.65,    273.65,  273.65,  273.65,
  273.8,     273.8,   273.8,   273.8,
  274.1,     274.1,   274.1,   274.1,
  274.55,    274.55,  274.55,  274.55,
  275,       275,     275,     275,
  275.5,     275.5,   275.5,   275.5,
  276,       276,     276,     276,
  276.5,     276.5,   276.5,   276.5,
  276.95,    276.95,  276.95,  276.95,
  277.35,    277.35,  277.35,  277.35,
  277.75,    277.75,  277.75,  277.75,
  278.05,    278.05,  278.05,  278.05,
  278.15,    278.15,  278.15,  278.15,
  278.25,    278.25,  278.25,  278.25,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.3,     278.3,   278.3,   278.3,
  278.2,     278.2,   278.2,   278.2,
  278.1,     278.1,   278.1,   278.1,
  278,       278,     278,     278,
  277.9,     277.9,   277.9,   277.9,
  277.8,     277.8,   277.8,   277.8,
  277.7,     277.7,   277.7,   277.7,
  277.65,    277.65,  277.65,  277.65,
  277.6,     277.6,   277.6,   277.6,
  277.45,    277.45,  277.45,  277.45,
  277.25,    277.25,  277.25,  277.25,
  277.1,     277.1,   277.1,   277.1,
  277,       277,     277,     277,
  276.9,     276.9,   276.9,   276.9,
  276.85,    276.85,  276.85,  276.85,
  276.85,    276.85,  276.85,  276.85,
  276.8,     276.8,   276.8,   276.8,
  276.8,     276.8,   276.8,   276.8,
  276.9,     276.9,   276.9,   276.9,
  276.95,    276.95,  276.95,  276.95,
  276.95,    276.95,  276.95,  276.95,
  276.9,     276.9,   276.9,   276.9,
  276.85,    276.85,  276.85,  276.85,
  276.85,    276.85,  276.85,  276.85,
  276.8,     276.8,   276.8,   276.8,
  276.7,     276.7,   276.7,   276.7,
  276.7,     276.7,   276.7,   276.7,
  276.75,    276.75,  276.75,  276.75,
  276.8,     276.8,   276.8,   276.8,
  276.9,     276.9,   276.9,   276.9,
  276.95,    276.95,  276.95,  276.95,
  276.85,    276.85,  276.85,  276.85,
  276.7,     276.7,   276.7,   276.7,
  276.8,     276.8,   276.8,   276.8,
  277.1,     277.1,   277.1,   277.1,
  277.35,    277.35,  277.35,  277.35,
  277.55,    277.55,  277.55,  277.55,
  277.75,    277.75,  277.75,  277.75,
  277.9,     277.9,   277.9,   277.9,
  277.85,    277.85,  277.85,  277.85,
  277.6,     277.6,   277.6,   277.6,
  277.35,    277.35,  277.35,  277.35,
  277.2,     277.2,   277.2,   277.2,
  277.1,     277.1,   277.1,   277.1,
  277,       277,     277,     277,
  277,       277,     277,     277,
  277.05,    277.05,  277.05,  277.05,
  277.1,     277.1,   277.1,   277.1,
  277.1,     277.1,   277.1,   277.1,
  277.1,     277.1,   277.1,   277.1,
  277.15,    277.15,  277.15,  277.15,
  277.15,    277.15,  277.15,  277.15,
  277.15,    277.15,  277.15,  277.15,
  277.15,    277.15,  277.15,  277.15,
  277.1,     277.1,   277.1,   277.1,
  277,       277,     277,     277,
  276.9,     276.9,   276.9,   276.9,
  276.85,    276.85,  276.85,  276.85,
  276.8,     276.8,   276.8,   276.8,
  276.75,    276.75,  276.75,  276.75,
  276.8,     276.8,   276.8,   276.8,
  276.85,    276.85,  276.85,  276.85,
  276.85,    276.85,  276.85,  276.85,
  276.9,     276.9,   276.9,   276.9,
  276.95,    276.95,  276.95,  276.95,
  277,       277,     277,     277,
  277.05,    277.05,  277.05,  277.05,
  277.05,    277.05,  277.05,  277.05,
  277.1,     277.1,   277.1,   277.1,
  277.15,    277.15,  277.15,  277.15,
  277.2,     277.2,   277.2,   277.2,
  277.25,    277.25,  277.25,  277.25,
  277.3,     277.3,   277.3,   277.3,
  277.35,    277.35,  277.35,  277.35,
  277.4,     277.4,   277.4,   277.4,
  277.45,    277.45,  277.45,  277.45,
  277.5,     277.5,   277.5,   277.5,
  277.65,    277.65,  277.65,  277.65,
  277.85,    277.85,  277.85,  277.85,
  278.05,    278.05,  278.05,  278.05,
  278.2,     278.2,   278.2,   278.2,
  278.3,     278.3,   278.3,   278.3,
  278.35,    278.35,  278.35,  278.35,
  278.45,    278.45,  278.45,  278.45,
  278.65,    278.65,  278.65,  278.65,
  278.9,     278.9,   278.9,   278.9,
  279.15,    279.15,  279.15,  279.15,
  279.4,     279.4,   279.4,   279.4,
  279.55,    279.55,  279.55,  279.55,
  279.55,    279.55,  279.55,  279.55,
  279.5,     279.5,   279.5,   279.5,
  279.35,    279.35,  279.35,  279.35,
  279.25,    279.25,  279.25,  279.25,
  279.25,    279.25,  279.25,  279.25,
  279.3,     279.3,   279.3,   279.3,
  279.45,    279.45,  279.45,  279.45,
  279.65,    279.65,  279.65,  279.65,
  279.8,     279.8,   279.8,   279.8,
  279.9,     279.9,   279.9,   279.9,
  280.1,     280.1,   280.1,   280.1,
  280.3,     280.3,   280.3,   280.3,
  280.5,     280.5,   280.5,   280.5,
  280.8,     280.8,   280.8,   280.8,
  281.05,    281.05,  281.05,  281.05,
  281.2,     281.2,   281.2,   281.2,
  281.3,     281.3,   281.3,   281.3,
  281.35,    281.35,  281.35,  281.35,
  281.35,    281.35,  281.35,  281.35,
  281.2,     281.2,   281.2,   281.2,
  281,       281,     281,     281,
  281,       281,     281,     281,
  281.05,    281.05,  281.05,  281.05,
  281.05,    281.05,  281.05,  281.05,
  281.1,     281.1,   281.1,   281.1,
  281.2,     281.2,   281.2,   281.2,
  281.25,    281.25,  281.25,  281.25,
  281.25,    281.25,  281.25,  281.25,
  281.25,    281.25,  281.25,  281.25,
  281.35,    281.35,  281.35,  281.35,
  281.5,     281.5,   281.5,   281.5,
  281.6,     281.6,   281.6,   281.6,
  281.65,    281.65,  281.65,  281.65,
  281.65,    281.65,  281.65,  281.65,
  281.6,     281.6,   281.6,   281.6,
  281.55,    281.55,  281.55,  281.55,
  281.55,    281.55,  281.55,  281.55,
  281.6,     281.6,   281.6,   281.6,
  281.7,     281.7,   281.7,   281.7,
  281.8,     281.8,   281.8,   281.8,
  281.95,    281.95,  281.95,  281.95,
  282.2,     282.2,   282.2,   282.2,
  282.45,    282.45,  282.45,  282.45,
  282.6,     282.6,   282.6,   282.6,
  282.85,    282.85,  282.85,  282.85,
  283.05,    283.05,  283.05,  283.05,
  283.15,    283.15,  283.15,  283.15,
  283.4,     283.4,   283.4,   283.4,
  283.55,    283.55,  283.55,  283.55,
  283.55,    283.55,  283.55,  283.55,
  283.55,    283.55,  283.55,  283.55,
  283.5,     283.5,   283.5,   283.5,
  283.25,    283.25,  283.25,  283.25,
  283.05,    283.05,  283.05,  283.05,
  283.05,    283.05,  283.05,  283.05,
  283.05,    283.05,  283.05,  283.05,
  283,       283,     283,     283,
  282.95,    282.95,  282.95,  282.95,
  282.85,    282.85,  282.85,  282.85,
  282.75,    282.75,  282.75,  282.75,
  282.7,     282.7,   282.7,   282.7,
  282.55,    282.55,  282.55,  282.55,
  282.35,    282.35,  282.35,  282.35,
  282.25,    282.25,  282.25,  282.25,
  282.2,     282.2,   282.2,   282.2,
  282.1,     282.1,   282.1,   282.1,
  281.9,     281.9,   281.9,   281.9,
  281.7,     281.7,   281.7,   281.7,
  281.55,    281.55,  281.55,  281.55,
  281.4,     281.4,   281.4,   281.4,
  281.45,    281.45,  281.45,  281.45,
  281.5,     281.5,   281.5,   281.5,
  281.5,     281.5,   281.5,   281.5,
  281.55,    281.55,  281.55,  281.55,
  281.55,    281.55,  281.55,  281.55,
  281.55,    281.55,  281.55,  281.55,
  281.5,     281.5,   281.5,   281.5,
  281.4,     281.4,   281.4,   281.4,
  281.25,    281.25,  281.25,  281.25,
  281.15,    281.15,  281.15,  281.15,
  281.15,    281.15,  281.15,  281.15,
  281.15,    281.15,  281.15,  281.15,
  281.2,     281.2,   281.2,   281.2,
  281.25,    281.25,  281.25,  281.25,
  281.2,     281.2,   281.2,   281.2,
  281.15,    281.15,  281.15,  281.15,
  281.2,     281.2,   281.2,   281.2,
  281.25,    281.25,  281.25,  281.25,
  281.2,     281.2,   281.2,   281.2,
  281.2,     281.2,   281.2,   281.2,
  281.25,    281.25,  281.25,  281.25,
  281.2,     281.2,   281.2,   281.2,
  281.2,     281.2,   281.2,   281.2,
  281.25,    281.25,  281.25,  281.25,
  281.3,     281.3,   281.3,   281.3,
  281.3,     281.3,   281.3,   281.3,
  281.25,    281.25,  281.25,  281.25,
  281.2,     281.2,   281.2,   281.2,
  281.1,     281.1,   281.1,   281.1,
  281.1,     281.1,   281.1,   281.1,
  281.15,    281.15,  281.15,  281.15,
  281.1,     281.1,   281.1,   281.1,
  281.05,    281.05,  281.05,  281.05,
  281,       281,     281,     281,
  280.95,    280.95,  280.95,  280.95,
  280.9,     280.9,   280.9,   280.9,
  280.8,     280.8,   280.8,   280.8,
  280.55,    280.55,  280.55,  280.55,
  279.9,     279.9,   279.9,   279.9,
  279.05,    279.05,  279.05,  279.05,
  278.45,    278.45,  278.45,  278.45,
  278.15,    278.15,  278.15,  278.15,
  278,       278,     278,     278,
  277.95,    277.95,  277.95,  277.95,
  277.95,    277.95,  277.95,  277.95,
  277.95,    277.95,  277.95,  277.95,
  277.95,    277.95,  277.95,  277.95,
  277.9,     277.9,   277.9,   277.9,
  277.65,    277.65,  277.65,  277.65,
  277.05,    277.05,  277.05,  277.05,
  276.4,     276.4,   276.4,   276.4,
  275.9,     275.9,   275.9,   275.9,
  275.45,    275.45,  275.45,  275.45,
  275.1,     275.1,   275.1,   275.1,
  274.8,     274.8,   274.8,   274.8,
  274.7,     274.7,   274.7,   274.7,
  274.7,     274.7,   274.7,   274.7,
  274.65,    274.65,  274.65,  274.65,
  274.55,    274.55,  274.55,  274.55,
  274.25,    274.25,  274.25,  274.25,
  274.2,     274.2,   274.2,   274.2,
  274.35,    274.35,  274.35,  274.35,
  274.25,    274.25,  274.25,  274.25,
  274.15,    274.15,  274.15,  274.15,
  273.8,     273.8,   273.8,   273.8,
  273.6,     273.6,   273.6,   273.6,
  274.15,    274.15,  274.15,  274.15,
  274.95,    274.95,  274.95,  274.95,
  275.9,     275.9,   275.9,   275.9,
  277.1,     277.1,   277.1,   277.1,
  278.25,    278.25,  278.25,  278.25,
  279.05,    279.05,  279.05,  279.05,
  279.5,     279.5,   279.5,   279.5,
  279.35,    279.35,  279.35,  279.35,
  279.25,    279.25,  279.25,  279.25,
  279.55,    279.55,  279.55,  279.55,
  279.25,    279.25,  279.25,  279.25,
  278.8,     278.8,   278.8,   278.8,
  278.55,    278.55,  278.55,  278.55,
  278.05,    278.05,  278.05,  278.05,
  277.55,    277.55,  277.55,  277.55,
  277,       277,     277,     277,
  276.35,    276.35,  276.35,  276.35,
  275.85,    275.85,  275.85,  275.85,
  275.35,    275.35,  275.35,  275.35,
  275.1,     275.1,   275.1,   275.1,
  274.9,     274.9,   274.9,   274.9,
  274.65,    274.65,  274.65,  274.65,
  274.7,     274.7,   274.7,   274.7,
  274.7,     274.7,   274.7,   274.7,
  274.8,     274.8,   274.8,   274.8,
  275,       275,     275,     275,
  275.05,    275.05,  275.05,  275.05,
  275,       275,     275,     275,
  275.05,    275.05,  275.05,  275.05,
  275.2,     275.2,   275.2,   275.2,
  275.35,    275.35,  275.35,  275.35,
  275.4,     275.4,   275.4,   275.4,
  275.3,     275.3,   275.3,   275.3,
  275.25,    275.25,  275.25,  275.25,
  275.25,    275.25,  275.25,  275.25,
  275.3,     275.3,   275.3,   275.3,
  275.35,    275.35,  275.35,  275.35,
  275.2,     275.2,   275.2,   275.2,
  274.85,    274.85,  274.85,  274.85,
  274.5,     274.5,   274.5,   274.5,
  274.15,    274.15,  274.15,  274.15,
  273.8,     273.8,   273.8,   273.8,
  273.6,     273.6,   273.6,   273.6,
  273.5,     273.5,   273.5,   273.5,
  273.45,    273.45,  273.45,  273.45,
  273.45,    273.45,  273.45,  273.45,
  273.45,    273.45,  273.45,  273.45,
  273.4,     273.4,   273.4,   273.4,
  273.4,     273.4,   273.4,   273.4,
  273.55,    273.55,  273.55,  273.55,
  273.9,     273.9,   273.9,   273.9,
  274.3,     274.3,   274.3,   274.3,
  274.6,     274.6,   274.6,   274.6,
  274.75,    274.75,  274.75,  274.75,
  274.85,    274.85,  274.85,  274.85,
  275.05,    275.05,  275.05,  275.05,
  275.15,    275.15,  275.15,  275.15,
  275.1,     275.1,   275.1,   275.1,
  275.05,    275.05,  275.05,  275.05,
  275,       275,     275,     275,
  274.85,    274.85,  274.85,  274.85,
  274.7,     274.7,   274.7,   274.7,
  274.65,    274.65,  274.65,  274.65,
  274.65,    274.65,  274.65,  274.65,
  274.6,     274.6,   274.6,   274.6,
  274.5,     274.5,   274.5,   274.5,
  274.4,     274.4,   274.4,   274.4,
  274.25,    274.25,  274.25,  274.25,
  274.05,    274.05,  274.05,  274.05,
  273.9,     273.9,   273.9,   273.9,
  273.8,     273.8,   273.8,   273.8,
  273.55,    273.55,  273.55,  273.55,
  273.35,    273.35,  273.35,  273.35,
  273.25,    273.25,  273.25,  273.25,
  273.2,     273.2,   273.2,   273.2,
  273.35,    273.35,  273.35,  273.35,
  273.5,     273.5,   273.5,   273.5,
  273.55,    273.55,  273.55,  273.55,
  273.55,    273.55,  273.55,  273.55,
  273.5,     273.5,   273.5,   273.5,
  273.35,    273.35,  273.35,  273.35,
  273.35,    273.35,  273.35,  273.35,
  273.55,    273.55,  273.55,  273.55,
  273.65,    273.65,  273.65,  273.65,
  273.55,    273.55,  273.55,  273.55,
  273.35,    273.35,  273.35,  273.35,
  273.15,    273.15,  273.15,  273.15,
  272.9,     272.9,   272.9,   272.9,
  272.65,    272.65,  272.65,  272.65,
  272.35,    272.35,  272.35,  272.35,
  271.95,    271.95,  271.95,  271.95,
  271.65,    271.65,  271.65,  271.65,
  271.5,     271.5,   271.5,   271.5,
  271.5,     271.5,   271.5,   271.5,
  271.55,    271.55,  271.55,  271.55,
  271.6,     271.6,   271.6,   271.6,
  271.65,    271.65,  271.65,  271.65,
  271.85,    271.85,  271.85,  271.85,
  272.35,    272.35,  272.35,  272.35,
  273.05,    273.05,  273.05,  273.05,
  273.95,    273.95,  273.95,  273.95,
  275.15,    275.15,  275.15,  275.15,
  276.45,    276.45,  276.45,  276.45,
  277.2,     277.2,   277.2,   277.2,
  277.2,     277.2,   277.2,   277.2,
  276.9,     276.9,   276.9,   276.9,
  276.55,    276.55,  276.55,  276.55,
  276.15,    276.15,  276.15,  276.15,
  275.95,    275.95,  275.95,  275.95,
  275.8,     275.8,   275.8,   275.8,
  275.45,    275.45,  275.45,  275.45,
  275.15,    275.15,  275.15,  275.15,
  274.95,    274.95,  274.95,  274.95,
  274.85,    274.85,  274.85,  274.85,
  274.9,     274.9,   274.9,   274.9,
  275,       275,     275,     275,
  275.05,    275.05,  275.05,  275.05,
  274.95,    274.95,  274.95,  274.95,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.9,     274.9,   274.9,   274.9,
  274.85,    274.85,  274.85,  274.85,
  274.5,     274.5,   274.5,   274.5,
  274,       274,     274,     274,
  273.55,    273.55,  273.55,  273.55,
  273.25,    273.25,  273.25,  273.25,
  273.2,     273.2,   273.2,   273.2,
  273.35,    273.35,  273.35,  273.35,
  273.5,     273.5,   273.5,   273.5,
  273.6,     273.6,   273.6,   273.6,
  273.75,    273.75,  273.75,  273.75,
  274,       274,     274,     274,
  274.25,    274.25,  274.25,  274.25,
  274.4,     274.4,   274.4,   274.4,
  274.55,    274.55,  274.55,  274.55,
  274.65,    274.65,  274.65,  274.65,
  274.7,     274.7,   274.7,   274.7,
  274.7,     274.7,   274.7,   274.7,
  274.6,     274.6,   274.6,   274.6,
  274.65,    274.65,  274.65,  274.65,
  274.9,     274.9,   274.9,   274.9,
  275.2,     275.2,   275.2,   275.2,
  275.4,     275.4,   275.4,   275.4,
  275.45,    275.45,  275.45,  275.45,
  275.45,    275.45,  275.45,  275.45,
  275.4,     275.4,   275.4,   275.4,
  275.3,     275.3,   275.3,   275.3,
  275.25,    275.25,  275.25,  275.25,
  275.25,    275.25,  275.25,  275.25,
  275.2,     275.2,   275.2,   275.2,
  275.05,    275.05,  275.05,  275.05,
  274.95,    274.95,  274.95,  274.95,
  274.85,    274.85,  274.85,  274.85,
  274.55,    274.55,  274.55,  274.55,
  274.15,    274.15,  274.15,  274.15,
  273.65,    273.65,  273.65,  273.65,
  272.95,    272.95,  272.95,  272.95,
  272.4,     272.4,   272.4,   272.4,
  272.2,     272.2,   272.2,   272.2,
  272.2,     272.2,   272.2,   272.2,
  271.85,    271.85,  271.85,  271.85,
  271.4,     271.4,   271.4,   271.4,
  271.4,     271.4,   271.4,   271.4,
  271.3,     271.3,   271.3,   271.3,
  271.05,    271.05,  271.05,  271.05,
  270.65,    270.65,  270.65,  270.65,
  270,       270,     270,     270,
  270.2,     270.2,   270.2,   270.2,
  270.2,     270.2,   270.2,   270.2,
  269.3,     269.3,   269.3,   269.3,
  268.85,    268.85,  268.85,  268.85,
  268.95,    268.95,  268.95,  268.95,
  269.15,    269.15,  269.15,  269.15,
  269.35,    269.35,  269.35,  269.35,
  269.65,    269.65,  269.65,  269.65,
  269.85,    269.85,  269.85,  269.85,
  269.85,    269.85,  269.85,  269.85,
  269.95,    269.95,  269.95,  269.95,
  270.4,     270.4,   270.4,   270.4,
  270.9,     270.9,   270.9,   270.9,
  271.3,     271.3,   271.3,   271.3,
  271.55,    271.55,  271.55,  271.55,
  271.7,     271.7,   271.7,   271.7,
  271.7,     271.7,   271.7,   271.7,
  271.65,    271.65,  271.65,  271.65,
  271.8,     271.8,   271.8,   271.8,
  272.1,     272.1,   272.1,   272.1,
  272.5,     272.5,   272.5,   272.5,
  272.95,    272.95,  272.95,  272.95,
  273.3,     273.3,   273.3,   273.3,
  273.75,    273.75,  273.75,  273.75,
  274.25,    274.25,  274.25,  274.25,
  274.6,     274.6,   274.6,   274.6,
  274.85,    274.85,  274.85,  274.85,
  275.45,    275.45,  275.45,  275.45,
  276.1,     276.1,   276.1,   276.1,
  276.3,     276.3,   276.3,   276.3,
  276.4,     276.4,   276.4,   276.4,
  276.3,     276.3,   276.3,   276.3,
  276.1,     276.1,   276.1,   276.1,
  276.05,    276.05,  276.05,  276.05,
  275.95,    275.95,  275.95,  275.95,
  275.75,    275.75,  275.75,  275.75,
  275.55,    275.55,  275.55,  275.55,
  275.45,    275.45,  275.45,  275.45,
  275.3,     275.3,   275.3,   275.3,
  274.8,     274.8,   274.8,   274.8,
  274.35,    274.35,  274.35,  274.35,
  274.25,    274.25,  274.25,  274.25,
  274.3,     274.3,   274.3,   274.3,
  274.2,     274.2,   274.2,   274.2,
  273.95,    273.95,  273.95,  273.95,
  273.8,     273.8,   273.8,   273.8,
  273.75,    273.75,  273.75,  273.75,
  273.75,    273.75,  273.75,  273.75,
  273.7,     273.7,   273.7,   273.7,
  273.7,     273.7,   273.7,   273.7,
  273.85,    273.85,  273.85,  273.85,
  273.95,    273.95,  273.95,  273.95,
  274,       274,     274,     274,
  274.15,    274.15,  274.15,  274.15,
  274.25,    274.25,  274.25,  274.25,
  274.15,    274.15,  274.15,  274.15,
  274.1,     274.1,   274.1,   274.1,
  274.15,    274.15,  274.15,  274.15,
  274.25,    274.25,  274.25,  274.25,
  274.45,    274.45,  274.45,  274.45,
  274.55,    274.55,  274.55,  274.55,
  274.6,     274.6,   274.6,   274.6,
  274.7,     274.7,   274.7,   274.7,
  274.8,     274.8,   274.8,   274.8,
  274.85,    274.85,  274.85,  274.85,
  274.9,     274.9,   274.9,   274.9,
  274.95,    274.95,  274.95,  274.95,
  275,       275,     275,     275,
  275.15,    275.15,  275.15,  275.15,
  275.15,    275.15,  275.15,  275.15,
  274.9,     274.9,   274.9,   274.9,
  274.9,     274.9,   274.9,   274.9,
  275,       275,     275,     275,
  274.85,    274.85,  274.85,  274.85,
  274.75,    274.75,  274.75,  274.75,
  274.75,    274.75,  274.75,  274.75,
  274.85,    274.85,  274.85,  274.85,
  275,       275,     275,     275,
  275.25,    275.25,  275.25,  275.25,
  275.7,     275.7,   275.7,   275.7,
  276,       276,     276,     276,
  276.15,    276.15,  276.15,  276.15,
  276.25,    276.25,  276.25,  276.25,
  276.3,     276.3,   276.3,   276.3,
  276.35,    276.35,  276.35,  276.35,
  276.5,     276.5,   276.5,   276.5,
  276.85,    276.85,  276.85,  276.85,
  277.2,     277.2,   277.2,   277.2,
  277.5,     277.5,   277.5,   277.5,
  277.7,     277.7,   277.7,   277.7,
  277.85,    277.85,  277.85,  277.85,
  278,       278,     278,     278,
  278.1,     278.1,   278.1,   278.1,
  278.2,     278.2,   278.2,   278.2,
  278.25,    278.25,  278.25,  278.25,
  278.25,    278.25,  278.25,  278.25,
  278.3,     278.3,   278.3,   278.3,
  278.3,     278.3,   278.3,   278.3,
  278.25,    278.25,  278.25,  278.25,
  278.3,     278.3,   278.3,   278.3,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.4,     278.4,   278.4,   278.4,
  278.35,    278.35,  278.35,  278.35,
  278,       278,     278,     278,
  277.3,     277.3,   277.3,   277.3,
  276.55,    276.55,  276.55,  276.55,
  276.15,    276.15,  276.15,  276.15,
  276.1,     276.1,   276.1,   276.1,
  276.2,     276.2,   276.2,   276.2,
  276.25,    276.25,  276.25,  276.25,
  276.25,    276.25,  276.25,  276.25,
  276.25,    276.25,  276.25,  276.25,
  276.25,    276.25,  276.25,  276.25,
  276.2,     276.2,   276.2,   276.2,
  276.05,    276.05,  276.05,  276.05,
  275.7,     275.7,   275.7,   275.7,
  275.2,     275.2,   275.2,   275.2,
  274.7,     274.7,   274.7,   274.7,
  274.4,     274.4,   274.4,   274.4,
  274.4,     274.4,   274.4,   274.4,
  274.55,    274.55,  274.55,  274.55,
  274.75,    274.75,  274.75,  274.75,
  275,       275,     275,     275,
  275.3,     275.3,   275.3,   275.3,
  275.5,     275.5,   275.5,   275.5,
  275.7,     275.7,   275.7,   275.7,
  275.95,    275.95,  275.95,  275.95,
  276.05,    276.05,  276.05,  276.05,
  275.9,     275.9,   275.9,   275.9,
  275.7,     275.7,   275.7,   275.7,
  275.6,     275.6,   275.6,   275.6,
  275.45,    275.45,  275.45,  275.45,
  275.25,    275.25,  275.25,  275.25,
  275.2,     275.2,   275.2,   275.2,
  275.3,     275.3,   275.3,   275.3,
  275.45,    275.45,  275.45,  275.45,
  275.65,    275.65,  275.65,  275.65,
  275.7,     275.7,   275.7,   275.7,
  275.35,    275.35,  275.35,  275.35,
  274.95,    274.95,  274.95,  274.95,
  274.85,    274.85,  274.85,  274.85,
  274.9,     274.9,   274.9,   274.9,
  275.15,    275.15,  275.15,  275.15,
  275.3,     275.3,   275.3,   275.3,
  275.25,    275.25,  275.25,  275.25,
  275.2,     275.2,   275.2,   275.2,
  275.25,    275.25,  275.25,  275.25,
  275.5,     275.5,   275.5,   275.5,
  275.65,    275.65,  275.65,  275.65,
  275.65,    275.65,  275.65,  275.65,
  275.75,    275.75,  275.75,  275.75,
  276.05,    276.05,  276.05,  276.05,
  276.4,     276.4,   276.4,   276.4,
  276.65,    276.65,  276.65,  276.65,
  276.75,    276.75,  276.75,  276.75,
  276.7,     276.7,   276.7,   276.7,
  276.65,    276.65,  276.65,  276.65,
  276.4,     276.4,   276.4,   276.4,
  276.25,    276.25,  276.25,  276.25,
  276.45,    276.45,  276.45,  276.45,
  276.8,     276.8,   276.8,   276.8,
  277.2,     277.2,   277.2,   277.2,
  277.2,     277.2,   277.2,   277.2,
  276.95,    276.95,  276.95,  276.95,
  276.95,    276.95,  276.95,  276.95,
  277.25,    277.25,  277.25,  277.25,
  277.6,     277.6,   277.6,   277.6,
  277.9,     277.9,   277.9,   277.9,
  278,       278,     278,     278,
  277.95,    277.95,  277.95,  277.95,
  278.05,    278.05,  278.05,  278.05,
  278.25,    278.25,  278.25,  278.25,
  278.4,     278.4,   278.4,   278.4,
  278.5,     278.5,   278.5,   278.5,
  278.6,     278.6,   278.6,   278.6,
  278.8,     278.8,   278.8,   278.8,
  279.2,     279.2,   279.2,   279.2,
  279.55,    279.55,  279.55,  279.55,
  279.8,     279.8,   279.8,   279.8,
  280.1,     280.1,   280.1,   280.1,
  280.25,    280.25,  280.25,  280.25,
  280.25,    280.25,  280.25,  280.25,
  280.05,    280.05,  280.05,  280.05,
  279.95,    279.95,  279.95,  279.95,
  280.25,    280.25,  280.25,  280.25,
  280.7,     280.7,   280.7,   280.7,
  281,       281,     281,     281,
  281,       281,     281,     281,
  280.85,    280.85,  280.85,  280.85,
  280.75,    280.75,  280.75,  280.75,
  280.85,    280.85,  280.85,  280.85,
  281,       281,     281,     281,
  281.1,     281.1,   281.1,   281.1,
  281.25,    281.25,  281.25,  281.25,
  281.4,     281.4,   281.4,   281.4,
  281.55,    281.55,  281.55,  281.55,
  281.65,    281.65,  281.65,  281.65,
  281.65,    281.65,  281.65,  281.65,
  281.7,     281.7,   281.7,   281.7,
  281.8,     281.8,   281.8,   281.8,
  281.75,    281.75,  281.75,  281.75,
  281.6,     281.6,   281.6,   281.6,
  281.6,     281.6,   281.6,   281.6,
  281.7,     281.7,   281.7,   281.7,
  281.8,     281.8,   281.8,   281.8,
  281.8,     281.8,   281.8,   281.8,
  281.7,     281.7,   281.7,   281.7,
  281.65,    281.65,  281.65,  281.65,
  281.6,     281.6,   281.6,   281.6,
  281.45,    281.45,  281.45,  281.45,
  281.3,     281.3,   281.3,   281.3,
  281.3,     281.3,   281.3,   281.3,
  281.4,     281.4,   281.4,   281.4,
  281.6,     281.6,   281.6,   281.6,
  281.85,    281.85,  281.85,  281.85,
  282,       282,     282,     282,
  282.25,    282.25,  282.25,  282.25,
  282.5,     282.5,   282.5,   282.5,
  282.65,    282.65,  282.65,  282.65,
  282.75,    282.75,  282.75,  282.75,
  282.75,    282.75,  282.75,  282.75,
  282.75,    282.75,  282.75,  282.75,
  282.7,     282.7,   282.7,   282.7,
  282.6,     282.6,   282.6,   282.6,
  282.4,     282.4,   282.4,   282.4,
  282.2,     282.2,   282.2,   282.2,
  282.1,     282.1,   282.1,   282.1,
  282.1,     282.1,   282.1,   282.1,
  282.15,    282.15,  282.15,  282.15,
  282.05,    282.05,  282.05,  282.05,
  281.75,    281.75,  281.75,  281.75,
  281.35,    281.35,  281.35,  281.35,
  281.2,     281.2,   281.2,   281.2,
  281.35,    281.35,  281.35,  281.35,
  281.5,     281.5,   281.5,   281.5,
  281.65,    281.65,  281.65,  281.65,
  281.8,     281.8,   281.8,   281.8,
  281.95,    281.95,  281.95,  281.95,
  282.15,    282.15,  282.15,  282.15,
  282.3,     282.3,   282.3,   282.3,
  282.4,     282.4,   282.4,   282.4,
  282.45,    282.45,  282.45,  282.45,
  282.45,    282.45,  282.45,  282.45,
  282.5,     282.5,   282.5,   282.5,
  282.6,     282.6,   282.6,   282.6,
  282.8,     282.8,   282.8,   282.8,
  283,       283,     283,     283,
  283.15,    283.15,  283.15,  283.15,
  283.3,     283.3,   283.3,   283.3,
  283.4,     283.4,   283.4,   283.4,
  283.45,    283.45,  283.45,  283.45,
  283.45,    283.45,  283.45,  283.45,
  283.4,     283.4,   283.4,   283.4,
  283.4,     283.4,   283.4,   283.4,
  283.45,    283.45,  283.45,  283.45,
  283.4,     283.4,   283.4,   283.4,
  283.35,    283.35,  283.35,  283.35,
  283.45,    283.45,  283.45,  283.45,
  283.65,    283.65,  283.65,  283.65,
  283.7,     283.7,   283.7,   283.7,
  283.65,    283.65,  283.65,  283.65,
  283.45,    283.45,  283.45,  283.45,
  283.15,    283.15,  283.15,  283.15,
  283,       283,     283,     283,
  282.95,    282.95,  282.95,  282.95,
  283,       283,     283,     283,
  283.15,    283.15,  283.15,  283.15,
  283.35,    283.35,  283.35,  283.35,
  283.6,     283.6,   283.6,   283.6,
  283.85,    283.85,  283.85,  283.85,
  284.05,    284.05,  284.05,  284.05,
  284.3,     284.3,   284.3,   284.3,
  284.65,    284.65,  284.65,  284.65,
  284.95,    284.95,  284.95,  284.95,
  285.15,    285.15,  285.15,  285.15,
  285.25,    285.25,  285.25,  285.25,
  285.1,     285.1,   285.1,   285.1,
  284.75,    284.75,  284.75,  284.75,
  284.45,    284.45,  284.45,  284.45,
  284.35,    284.35,  284.35,  284.35,
  284.45,    284.45,  284.45,  284.45,
  284.5,     284.5,   284.5,   284.5,
  284.45,    284.45,  284.45,  284.45,
  284.45,    284.45,  284.45,  284.45,
  284.45,    284.45,  284.45,  284.45,
  284.55,    284.55,  284.55,  284.55,
  284.7,     284.7,   284.7,   284.7,
  284.7,     284.7,   284.7,   284.7,
  284.55,    284.55,  284.55,  284.55,
  284.4,     284.4,   284.4,   284.4,
  284.2,     284.2,   284.2,   284.2,
  284,       284,     284,     284,
  283.95,    283.95,  283.95,  283.95,
  283.9,     283.9,   283.9,   283.9,
  283.8,     283.8,   283.8,   283.8,
  283.7,     283.7,   283.7,   283.7,
  283.45,    283.45,  283.45,  283.45,
  283.25,    283.25,  283.25,  283.25,
  283.3,     283.3,   283.3,   283.3,
  283.3,     283.3,   283.3,   283.3,
  283.35,    283.35,  283.35,  283.35,
  283.45,    283.45,  283.45,  283.45,
  283.5,     283.5,   283.5,   283.5,
  283.6,     283.6,   283.6,   283.6,
  283.65,    283.65,  283.65,  283.65,
  283.5,     283.5,   283.5,   283.5,
  283.25,    283.25,  283.25,  283.25,
  283.15,    283.15,  283.15,  283.15,
  283.1,     283.1,   283.1,   283.1,
  283.1,     283.1,   283.1,   283.1,
  283.35,    283.35,  283.35,  283.35,
  283.75,    283.75,  283.75,  283.75,
  284.25,    284.25,  284.25,  284.25,
  284.8,     284.8,   284.8,   284.8,
  285.15,    285.15,  285.15,  285.15,
  285.3,     285.3,   285.3,   285.3,
  285.45,    285.45,  285.45,  285.45,
  285.55,    285.55,  285.55,  285.55,
  285.5,     285.5,   285.5,   285.5,
  285.35,    285.35,  285.35,  285.35,
  285.2,     285.2,   285.2,   285.2,
  285.15,    285.15,  285.15,  285.15,
  285.1,     285.1,   285.1,   285.1,
  284.95,    284.95,  284.95,  284.95,
  284.75,    284.75,  284.75,  284.75,
  284.65,    284.65,  284.65,  284.65,
  284.65,    284.65,  284.65,  284.65,
  284.55,    284.55,  284.55,  284.55,
  284.3,     284.3,   284.3,   284.3,
  283.95,    283.95,  283.95,  283.95,
  283.65,    283.65,  283.65,  283.65,
  283.65,    283.65,  283.65,  283.65,
  283.7,     283.7,   283.7,   283.7,
  283.6,     283.6,   283.6,   283.6,
  283.55,    283.55,  283.55,  283.55,
  283.5,     283.5,   283.5,   283.5,
  283.2,     283.2,   283.2,   283.2,
  282.7,     282.7,   282.7,   282.7,
  282.25,    282.25,  282.25,  282.25,
  281.95,    281.95,  281.95,  281.95,
  281.85,    281.85,  281.85,  281.85,
  281.85,    281.85,  281.85,  281.85,
  281.8,     281.8,   281.8,   281.8,
  281.7,     281.7,   281.7,   281.7,
  281.5,     281.5,   281.5,   281.5,
  281.15,    281.15,  281.15,  281.15,
  280.9,     280.9,   280.9,   280.9,
  280.85,    280.85,  280.85,  280.85,
  281.05,    281.05,  281.05,  281.05,
  281.3,     281.3,   281.3,   281.3,
  281.4,     281.4,   281.4,   281.4,
  281.2,     281.2,   281.2,   281.2,
  280.9,     280.9,   280.9,   280.9,
  280.8,     280.8,   280.8,   280.8,
  280.55,    280.55,  280.55,  280.55,
  280.25,    280.25,  280.25,  280.25,
  280.15,    280.15,  280.15,  280.15,
  280.2,     280.2,   280.2,   280.2,
  280.4,     280.4,   280.4,   280.4,
  280.7,     280.7,   280.7,   280.7,
  280.75,    280.75,  280.75,  280.75,
  280.6,     280.6,   280.6,   280.6,
  280.6,     280.6,   280.6,   280.6,
  280.75,    280.75,  280.75,  280.75,
  280.9,     280.9,   280.9,   280.9,
  280.95,    280.95,  280.95,  280.95,
  281,       281,     281,     281,
  281,       281,     281,     281,
  280.8,     280.8,   280.8,   280.8,
  280.45,    280.45,  280.45,  280.45,
  280.15,    280.15,  280.15,  280.15,
  280.1,     280.1,   280.1,   280.1,
  280.15,    280.15,  280.15,  280.15,
  280.05,    280.05,  280.05,  280.05,
  279.85,    279.85,  279.85,  279.85,
  279.7,     279.7,   279.7,   279.7,
  279.65,    279.65,  279.65,  279.65,
  279.7,     279.7,   279.7,   279.7,
  279.7,     279.7,   279.7,   279.7,
  279.45,    279.45,  279.45,  279.45,
  279.05,    279.05,  279.05,  279.05,
  278.8,     278.8,   278.8,   278.8,
  279,       279,     279,     279,
  279.35,    279.35,  279.35,  279.35,
  279.3,     279.3,   279.3,   279.3,
  279.05,    279.05,  279.05,  279.05,
  278.7,     278.7,   278.7,   278.7,
  278.5,     278.5,   278.5,   278.5,
  278.55,    278.55,  278.55,  278.55,
  278.3,     278.3,   278.3,   278.3,
  277.6,     277.6,   277.6,   277.6,
  277.05,    277.05,  277.05,  277.05,
  276.9,     276.9,   276.9,   276.9,
  276.85,    276.85,  276.85,  276.85,
  276.75,    276.75,  276.75,  276.75,
  276.6,     276.6,   276.6,   276.6,
  276.7,     276.7,   276.7,   276.7,
  277,       277,     277,     277,
  277.3,     277.3,   277.3,   277.3,
  277.35,    277.35,  277.35,  277.35,
  277.1,     277.1,   277.1,   277.1,
  276.8,     276.8,   276.8,   276.8,
  276.65,    276.65,  276.65,  276.65,
  276.65,    276.65,  276.65,  276.65,
  276.95,    276.95,  276.95,  276.95,
  277.5,     277.5,   277.5,   277.5,
  278.4,     278.4,   278.4,   278.4,
  279.65,    279.65,  279.65,  279.65,
  280.6,     280.6,   280.6,   280.6,
  281.15,    281.15,  281.15,  281.15,
  281.35,    281.35,  281.35,  281.35,
  281.3,     281.3,   281.3,   281.3,
  281.25,    281.25,  281.25,  281.25,
  281.1,     281.1,   281.1,   281.1,
  280.7,     280.7,   280.7,   280.7,
  280.45,    280.45,  280.45,  280.45,
  280.5,     280.5,   280.5,   280.5,
  280.65,    280.65,  280.65,  280.65,
  280.75,    280.75,  280.75,  280.75,
  280.8,     280.8,   280.8,   280.8,
  280.85,    280.85,  280.85,  280.85,
  280.85,    280.85,  280.85,  280.85,
  280.8,     280.8,   280.8,   280.8,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.55,    280.55,  280.55,  280.55,
  280.35,    280.35,  280.35,  280.35,
  280.1,     280.1,   280.1,   280.1,
  279.85,    279.85,  279.85,  279.85,
  279.6,     279.6,   279.6,   279.6,
  279.45,    279.45,  279.45,  279.45,
  279.4,     279.4,   279.4,   279.4,
  279.25,    279.25,  279.25,  279.25,
  279.1,     279.1,   279.1,   279.1,
  278.9,     278.9,   278.9,   278.9,
  278.65,    278.65,  278.65,  278.65,
  278.55,    278.55,  278.55,  278.55,
  278.55,    278.55,  278.55,  278.55,
  278.6,     278.6,   278.6,   278.6,
  278.65,    278.65,  278.65,  278.65,
  278.5,     278.5,   278.5,   278.5,
  278.35,    278.35,  278.35,  278.35,
  278.2,     278.2,   278.2,   278.2,
  277.95,    277.95,  277.95,  277.95,
  277.65,    277.65,  277.65,  277.65,
  277.4,     277.4,   277.4,   277.4,
  277.25,    277.25,  277.25,  277.25,
  276.95,    276.95,  276.95,  276.95,
  276.75,    276.75,  276.75,  276.75,
  276.7,     276.7,   276.7,   276.7,
  276.55,    276.55,  276.55,  276.55,
  276.55,    276.55,  276.55,  276.55,
  276.85,    276.85,  276.85,  276.85,
  277.3,     277.3,   277.3,   277.3,
  278.05,    278.05,  278.05,  278.05,
  279,       279,     279,     279,
  279.75,    279.75,  279.75,  279.75,
  280.05,    280.05,  280.05,  280.05,
  280.2,     280.2,   280.2,   280.2,
  280.3,     280.3,   280.3,   280.3,
  280.15,    280.15,  280.15,  280.15,
  279.9,     279.9,   279.9,   279.9,
  279.65,    279.65,  279.65,  279.65,
  279.5,     279.5,   279.5,   279.5,
  278.9,     278.9,   278.9,   278.9,
  278.25,    278.25,  278.25,  278.25,
  277.95,    277.95,  277.95,  277.95,
  277.6,     277.6,   277.6,   277.6,
  277.35,    277.35,  277.35,  277.35,
  277.2,     277.2,   277.2,   277.2,
  277.15,    277.15,  277.15,  277.15,
  277.1,     277.1,   277.1,   277.1,
  277.1,     277.1,   277.1,   277.1,
  277.1,     277.1,   277.1,   277.1,
  277,       277,     277,     277,
  276.85,    276.85,  276.85,  276.85,
  276.55,    276.55,  276.55,  276.55,
  276.1,     276.1,   276.1,   276.1,
  275.65,    275.65,  275.65,  275.65,
  275.3,     275.3,   275.3,   275.3,
  275.05,    275.05,  275.05,  275.05,
  275.1,     275.1,   275.1,   275.1,
  275.4,     275.4,   275.4,   275.4,
  275.55,    275.55,  275.55,  275.55,
  275.25,    275.25,  275.25,  275.25,
  274.6,     274.6,   274.6,   274.6,
  274.1,     274.1,   274.1,   274.1,
  273.85,    273.85,  273.85,  273.85,
  273.9,     273.9,   273.9,   273.9,
  274.25,    274.25,  274.25,  274.25,
  274.65,    274.65,  274.65,  274.65,
  275.05,    275.05,  275.05,  275.05,
  275.4,     275.4,   275.4,   275.4,
  275.5,     275.5,   275.5,   275.5,
  275.45,    275.45,  275.45,  275.45,
  275.3,     275.3,   275.3,   275.3,
  274.95,    274.95,  274.95,  274.95,
  274.6,     274.6,   274.6,   274.6,
  274.5,     274.5,   274.5,   274.5,
  274.6,     274.6,   274.6,   274.6,
  274.75,    274.75,  274.75,  274.75,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.9,     274.9,   274.9,   274.9,
  275.05,    275.05,  275.05,  275.05,
  275.25,    275.25,  275.25,  275.25,
  275.4,     275.4,   275.4,   275.4,
  275.45,    275.45,  275.45,  275.45,
  275.45,    275.45,  275.45,  275.45,
  275.4,     275.4,   275.4,   275.4,
  275.3,     275.3,   275.3,   275.3,
  275.2,     275.2,   275.2,   275.2,
  275,       275,     275,     275,
  274.7,     274.7,   274.7,   274.7,
  274.5,     274.5,   274.5,   274.5,
  274.35,    274.35,  274.35,  274.35,
  274.15,    274.15,  274.15,  274.15,
  274,       274,     274,     274,
  273.9,     273.9,   273.9,   273.9,
  273.7,     273.7,   273.7,   273.7,
  273.4,     273.4,   273.4,   273.4,
  273.1,     273.1,   273.1,   273.1,
  272.9,     272.9,   272.9,   272.9,
  272.8,     272.8,   272.8,   272.8,
  272.55,    272.55,  272.55,  272.55,
  272.2,     272.2,   272.2,   272.2,
  271.9,     271.9,   271.9,   271.9,
  271.6,     271.6,   271.6,   271.6,
  271.3,     271.3,   271.3,   271.3,
  271.1,     271.1,   271.1,   271.1,
  271,       271,     271,     271,
  270.85,    270.85,  270.85,  270.85,
  270.75,    270.75,  270.75,  270.75,
  270.75,    270.75,  270.75,  270.75,
  270.8,     270.8,   270.8,   270.8,
  270.85,    270.85,  270.85,  270.85,
  270.85,    270.85,  270.85,  270.85,
  270.9,     270.9,   270.9,   270.9,
  271,       271,     271,     271,
  271.05,    271.05,  271.05,  271.05,
  271.05,    271.05,  271.05,  271.05,
  270.95,    270.95,  270.95,  270.95,
  270.8,     270.8,   270.8,   270.8,
  270.7,     270.7,   270.7,   270.7,
  270.65,    270.65,  270.65,  270.65,
  270.55,    270.55,  270.55,  270.55,
  270.35,    270.35,  270.35,  270.35,
  270.2,     270.2,   270.2,   270.2,
  270.15,    270.15,  270.15,  270.15,
  270.1,     270.1,   270.1,   270.1,
  269.75,    269.75,  269.75,  269.75,
  269.2,     269.2,   269.2,   269.2,
  268.9,     268.9,   268.9,   268.9,
  268.9,     268.9,   268.9,   268.9,
  269.1,     269.1,   269.1,   269.1,
  269.2,     269.2,   269.2,   269.2,
  269.05,    269.05,  269.05,  269.05,
  268.95,    268.95,  268.95,  268.95,
  268.95,    268.95,  268.95,  268.95,
  268.85,    268.85,  268.85,  268.85,
  268.65,    268.65,  268.65,  268.65,
  268.4,     268.4,   268.4,   268.4,
  268.1,     268.1,   268.1,   268.1,
  267.9,     267.9,   267.9,   267.9,
  267.7,     267.7,   267.7,   267.7,
  267.45,    267.45,  267.45,  267.45,
  267.35,    267.35,  267.35,  267.35,
  267.25,    267.25,  267.25,  267.25,
  267.1,     267.1,   267.1,   267.1,
  267,       267,     267,     267,
  266.9,     266.9,   266.9,   266.9,
  266.85,    266.85,  266.85,  266.85,
  266.85,    266.85,  266.85,  266.85,
  266.75,    266.75,  266.75,  266.75,
  266.55,    266.55,  266.55,  266.55,
  266.4,     266.4,   266.4,   266.4,
  266.35,    266.35,  266.35,  266.35,
  266.25,    266.25,  266.25,  266.25,
  266.1,     266.1,   266.1,   266.1,
  266,       266,     266,     266,
  265.9,     265.9,   265.9,   265.9,
  265.85,    265.85,  265.85,  265.85,
  265.85,    265.85,  265.85,  265.85,
  265.9,     265.9,   265.9,   265.9,
  265.95,    265.95,  265.95,  265.95,
  265.95,    265.95,  265.95,  265.95,
  265.9,     265.9,   265.9,   265.9,
  265.8,     265.8,   265.8,   265.8,
  265.75,    265.75,  265.75,  265.75,
  265.7,     265.7,   265.7,   265.7,
  265.65,    265.65,  265.65,  265.65,
  265.7,     265.7,   265.7,   265.7,
  265.75,    265.75,  265.75,  265.75,
  265.8,     265.8,   265.8,   265.8,
  265.85,    265.85,  265.85,  265.85,
  265.9,     265.9,   265.9,   265.9,
  266.1,     266.1,   266.1,   266.1,
  266.45,    266.45,  266.45,  266.45,
  266.85,    266.85,  266.85,  266.85,
  267.35,    267.35,  267.35,  267.35,
  267.9,     267.9,   267.9,   267.9,
  268.25,    268.25,  268.25,  268.25,
  268.55,    268.55,  268.55,  268.55,
  269,       269,     269,     269,
  269.5,     269.5,   269.5,   269.5,
  269.9,     269.9,   269.9,   269.9,
  270.2,     270.2,   270.2,   270.2,
  270.55,    270.55,  270.55,  270.55,
  270.8,     270.8,   270.8,   270.8,
  270.95,    270.95,  270.95,  270.95,
  271.05,    271.05,  271.05,  271.05,
  271.15,    271.15,  271.15,  271.15,
  271.3,     271.3,   271.3,   271.3,
  271.35,    271.35,  271.35,  271.35,
  271.35,    271.35,  271.35,  271.35,
  271.3,     271.3,   271.3,   271.3,
  271.25,    271.25,  271.25,  271.25,
  271.3,     271.3,   271.3,   271.3,
  271.35,    271.35,  271.35,  271.35,
  271.35,    271.35,  271.35,  271.35,
  271.4,     271.4,   271.4,   271.4,
  271.5,     271.5,   271.5,   271.5,
  271.55,    271.55,  271.55,  271.55,
  271.6,     271.6,   271.6,   271.6,
  271.7,     271.7,   271.7,   271.7,
  271.8,     271.8,   271.8,   271.8,
  271.95,    271.95,  271.95,  271.95,
  272.2,     272.2,   272.2,   272.2,
  272.55,    272.55,  272.55,  272.55,
  272.85,    272.85,  272.85,  272.85,
  273.05,    273.05,  273.05,  273.05,
  273.25,    273.25,  273.25,  273.25,
  273.4,     273.4,   273.4,   273.4,
  273.4,     273.4,   273.4,   273.4,
  273.35,    273.35,  273.35,  273.35,
  273.55,    273.55,  273.55,  273.55,
  274.05,    274.05,  274.05,  274.05,
  274.4,     274.4,   274.4,   274.4,
  274.4,     274.4,   274.4,   274.4,
  274.3,     274.3,   274.3,   274.3,
  274.35,    274.35,  274.35,  274.35,
  274.8,     274.8,   274.8,   274.8,
  274.85,    274.85,  274.85,  274.85,
  274.8,     274.8,   274.8,   274.8,
  275.45,    275.45,  275.45,  275.45,
  276.1,     276.1,   276.1,   276.1,
  276.6,     276.6,   276.6,   276.6,
  277.05,    277.05,  277.05,  277.05,
  277.6,     277.6,   277.6,   277.6,
  278,       278,     278,     278,
  278,       278,     278,     278,
  278.05,    278.05,  278.05,  278.05,
  278.15,    278.15,  278.15,  278.15,
  278.25,    278.25,  278.25,  278.25,
  278.4,     278.4,   278.4,   278.4,
  278.5,     278.5,   278.5,   278.5,
  278.8,     278.8,   278.8,   278.8,
  278.95,    278.95,  278.95,  278.95,
  278.45,    278.45,  278.45,  278.45,
  277.95,    277.95,  277.95,  277.95,
  277.9,     277.9,   277.9,   277.9,
  278.05,    278.05,  278.05,  278.05,
  278.3,     278.3,   278.3,   278.3,
  278.55,    278.55,  278.55,  278.55,
  278.7,     278.7,   278.7,   278.7,
  278.8,     278.8,   278.8,   278.8,
  278.65,    278.65,  278.65,  278.65,
  278.2,     278.2,   278.2,   278.2,
  278.05,    278.05,  278.05,  278.05,
  278,       278,     278,     278,
  277.75,    277.75,  277.75,  277.75,
  277.45,    277.45,  277.45,  277.45,
  277.25,    277.25,  277.25,  277.25,
  277.35,    277.35,  277.35,  277.35,
  277.45,    277.45,  277.45,  277.45,
  277.5,     277.5,   277.5,   277.5,
  277.6,     277.6,   277.6,   277.6,
  277.7,     277.7,   277.7,   277.7,
  277.5,     277.5,   277.5,   277.5,
  277.15,    277.15,  277.15,  277.15,
  277.05,    277.05,  277.05,  277.05,
  277.1,     277.1,   277.1,   277.1,
  277.2,     277.2,   277.2,   277.2,
  277.3,     277.3,   277.3,   277.3,
  277.45,    277.45,  277.45,  277.45,
  277.65,    277.65,  277.65,  277.65,
  277.85,    277.85,  277.85,  277.85,
  278,       278,     278,     278,
  278.15,    278.15,  278.15,  278.15,
  278.45,    278.45,  278.45,  278.45,
  278.85,    278.85,  278.85,  278.85,
  279.1,     279.1,   279.1,   279.1,
  279.2,     279.2,   279.2,   279.2,
  279.3,     279.3,   279.3,   279.3,
  279.4,     279.4,   279.4,   279.4,
  279.5,     279.5,   279.5,   279.5,
  279.65,    279.65,  279.65,  279.65,
  280.1,     280.1,   280.1,   280.1,
  280.8,     280.8,   280.8,   280.8,
  281.35,    281.35,  281.35,  281.35,
  281.6,     281.6,   281.6,   281.6,
  281.5,     281.5,   281.5,   281.5,
  281.4,     281.4,   281.4,   281.4,
  281.75,    281.75,  281.75,  281.75,
  282.2,     282.2,   282.2,   282.2,
  282.3,     282.3,   282.3,   282.3,
  282.2,     282.2,   282.2,   282.2,
  282.3,     282.3,   282.3,   282.3,
  282.45,    282.45,  282.45,  282.45,
  282.35,    282.35,  282.35,  282.35,
  282.1,     282.1,   282.1,   282.1,
  281.6,     281.6,   281.6,   281.6,
  280.9,     280.9,   280.9,   280.9,
  280.65,    280.65,  280.65,  280.65,
  280.8,     280.8,   280.8,   280.8,
  280.85,    280.85,  280.85,  280.85,
  280.8,     280.8,   280.8,   280.8,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.55,    280.55,  280.55,  280.55,
  280.2,     280.2,   280.2,   280.2,
  279.8,     279.8,   279.8,   279.8,
  279.5,     279.5,   279.5,   279.5,
  279.25,    279.25,  279.25,  279.25,
  278.95,    278.95,  278.95,  278.95,
  278.55,    278.55,  278.55,  278.55,
  278.15,    278.15,  278.15,  278.15,
  277.7,     277.7,   277.7,   277.7,
  277.25,    277.25,  277.25,  277.25,
  276.85,    276.85,  276.85,  276.85,
  276.55,    276.55,  276.55,  276.55,
  276.3,     276.3,   276.3,   276.3,
  276.05,    276.05,  276.05,  276.05,
  275.85,    275.85,  275.85,  275.85,
  275.75,    275.75,  275.75,  275.75,
  275.8,     275.8,   275.8,   275.8,
  275.75,    275.75,  275.75,  275.75,
  275.3,     275.3,   275.3,   275.3,
  274.75,    274.75,  274.75,  274.75,
  274.45,    274.45,  274.45,  274.45,
  274.4,     274.4,   274.4,   274.4,
  274.75,    274.75,  274.75,  274.75,
  275.25,    275.25,  275.25,  275.25,
  275.75,    275.75,  275.75,  275.75,
  276.15,    276.15,  276.15,  276.15,
  276.55,    276.55,  276.55,  276.55,
  277.2,     277.2,   277.2,   277.2,
  277.75,    277.75,  277.75,  277.75,
  278,       278,     278,     278,
  278.25,    278.25,  278.25,  278.25,
  278.55,    278.55,  278.55,  278.55,
  278.55,    278.55,  278.55,  278.55,
  278.25,    278.25,  278.25,  278.25,
  277.6,     277.6,   277.6,   277.6,
  276.75,    276.75,  276.75,  276.75,
  276.1,     276.1,   276.1,   276.1,
  275.7,     275.7,   275.7,   275.7,
  275.45,    275.45,  275.45,  275.45,
  275.3,     275.3,   275.3,   275.3,
  275.2,     275.2,   275.2,   275.2,
  275.25,    275.25,  275.25,  275.25,
  275.4,     275.4,   275.4,   275.4,
  275.45,    275.45,  275.45,  275.45,
  275.4,     275.4,   275.4,   275.4,
  275.4,     275.4,   275.4,   275.4,
  275.7,     275.7,   275.7,   275.7,
  276.1,     276.1,   276.1,   276.1,
  276.2,     276.2,   276.2,   276.2,
  276.3,     276.3,   276.3,   276.3,
  276.2,     276.2,   276.2,   276.2,
  275.8,     275.8,   275.8,   275.8,
  275.7,     275.7,   275.7,   275.7,
  275.7,     275.7,   275.7,   275.7,
  275.55,    275.55,  275.55,  275.55,
  275.35,    275.35,  275.35,  275.35,
  275.2,     275.2,   275.2,   275.2,
  275.15,    275.15,  275.15,  275.15,
  275.1,     275.1,   275.1,   275.1,
  274.95,    274.95,  274.95,  274.95,
  274.8,     274.8,   274.8,   274.8,
  274.7,     274.7,   274.7,   274.7,
  274.6,     274.6,   274.6,   274.6,
  274.5,     274.5,   274.5,   274.5,
  274.5,     274.5,   274.5,   274.5,
  274.6,     274.6,   274.6,   274.6,
  274.65,    274.65,  274.65,  274.65,
  274.7,     274.7,   274.7,   274.7,
  274.85,    274.85,  274.85,  274.85,
  275,       275,     275,     275,
  275.15,    275.15,  275.15,  275.15,
  275.35,    275.35,  275.35,  275.35,
  275.45,    275.45,  275.45,  275.45,
  275.5,     275.5,   275.5,   275.5,
  275.55,    275.55,  275.55,  275.55,
  275.55,    275.55,  275.55,  275.55,
  275.55,    275.55,  275.55,  275.55,
  275.55,    275.55,  275.55,  275.55,
  275.6,     275.6,   275.6,   275.6,
  275.65,    275.65,  275.65,  275.65,
  275.7,     275.7,   275.7,   275.7,
  275.75,    275.75,  275.75,  275.75,
  275.75,    275.75,  275.75,  275.75,
  275.75,    275.75,  275.75,  275.75,
  275.75,    275.75,  275.75,  275.75,
  275.7,     275.7,   275.7,   275.7,
  275.55,    275.55,  275.55,  275.55,
  275.45,    275.45,  275.45,  275.45,
  275.45,    275.45,  275.45,  275.45,
  275.45,    275.45,  275.45,  275.45,
  275.45,    275.45,  275.45,  275.45,
  275.5,     275.5,   275.5,   275.5,
  275.55,    275.55,  275.55,  275.55,
  275.6,     275.6,   275.6,   275.6,
  275.7,     275.7,   275.7,   275.7,
  275.75,    275.75,  275.75,  275.75,
  275.8,     275.8,   275.8,   275.8,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.8,     275.8,   275.8,   275.8,
  275.7,     275.7,   275.7,   275.7,
  275.6,     275.6,   275.6,   275.6,
  275.55,    275.55,  275.55,  275.55,
  275.5,     275.5,   275.5,   275.5,
  275.45,    275.45,  275.45,  275.45,
  275.35,    275.35,  275.35,  275.35,
  275.2,     275.2,   275.2,   275.2,
  275.05,    275.05,  275.05,  275.05,
  274.9,     274.9,   274.9,   274.9,
  274.8,     274.8,   274.8,   274.8,
  274.7,     274.7,   274.7,   274.7,
  274.6,     274.6,   274.6,   274.6,
  274.55,    274.55,  274.55,  274.55,
  274.5,     274.5,   274.5,   274.5,
  274.5,     274.5,   274.5,   274.5,
  274.55,    274.55,  274.55,  274.55,
  274.6,     274.6,   274.6,   274.6,
  274.7,     274.7,   274.7,   274.7,
  274.8,     274.8,   274.8,   274.8,
  274.9,     274.9,   274.9,   274.9,
  275,       275,     275,     275,
  275.1,     275.1,   275.1,   275.1,
  275.15,    275.15,  275.15,  275.15,
  275.2,     275.2,   275.2,   275.2,
  275.25,    275.25,  275.25,  275.25,
  275.25,    275.25,  275.25,  275.25,
  275.25,    275.25,  275.25,  275.25,
  275.25,    275.25,  275.25,  275.25,
  275.25,    275.25,  275.25,  275.25,
  275.2,     275.2,   275.2,   275.2,
  275.15,    275.15,  275.15,  275.15,
  275.15,    275.15,  275.15,  275.15,
  275.1,     275.1,   275.1,   275.1,
  275.05,    275.05,  275.05,  275.05,
  275.05,    275.05,  275.05,  275.05,
  275,       275,     275,     275,
  274.95,    274.95,  274.95,  274.95,
  275,       275,     275,     275,
  275,       275,     275,     275,
  274.95,    274.95,  274.95,  274.95,
  274.95,    274.95,  274.95,  274.95,
  274.95,    274.95,  274.95,  274.95,
  274.95,    274.95,  274.95,  274.95,
  274.95,    274.95,  274.95,  274.95,
  274.9,     274.9,   274.9,   274.9,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.85,    274.85,  274.85,  274.85,
  274.8,     274.8,   274.8,   274.8,
  274.75,    274.75,  274.75,  274.75,
  274.7,     274.7,   274.7,   274.7,
  274.65,    274.65,  274.65,  274.65,
  274.6,     274.6,   274.6,   274.6,
  274.55,    274.55,  274.55,  274.55,
  274.5,     274.5,   274.5,   274.5,
  274.45,    274.45,  274.45,  274.45,
  274.45,    274.45,  274.45,  274.45,
  274.5,     274.5,   274.5,   274.5,
  274.6,     274.6,   274.6,   274.6,
  274.65,    274.65,  274.65,  274.65,
  274.7,     274.7,   274.7,   274.7,
  274.8,     274.8,   274.8,   274.8,
  274.9,     274.9,   274.9,   274.9,
  275,       275,     275,     275,
  275.2,     275.2,   275.2,   275.2,
  275.4,     275.4,   275.4,   275.4,
  275.55,    275.55,  275.55,  275.55,
  275.7,     275.7,   275.7,   275.7,
  275.75,    275.75,  275.75,  275.75,
  275.75,    275.75,  275.75,  275.75,
  275.8,     275.8,   275.8,   275.8,
  275.8,     275.8,   275.8,   275.8,
  275.8,     275.8,   275.8,   275.8,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.85,    275.85,  275.85,  275.85,
  275.9,     275.9,   275.9,   275.9,
  276.05,    276.05,  276.05,  276.05,
  276.25,    276.25,  276.25,  276.25,
  276.5,     276.5,   276.5,   276.5,
  276.85,    276.85,  276.85,  276.85,
  277.15,    277.15,  277.15,  277.15,
  277.4,     277.4,   277.4,   277.4,
  277.65,    277.65,  277.65,  277.65,
  277.85,    277.85,  277.85,  277.85,
  278,       278,     278,     278,
  278.1,     278.1,   278.1,   278.1,
  278.2,     278.2,   278.2,   278.2,
  278.3,     278.3,   278.3,   278.3,
  278.4,     278.4,   278.4,   278.4,
  278.55,    278.55,  278.55,  278.55,
  278.7,     278.7,   278.7,   278.7,
  278.8,     278.8,   278.8,   278.8,
  278.85,    278.85,  278.85,  278.85,
  278.9,     278.9,   278.9,   278.9,
  279,       279,     279,     279,
  279.1,     279.1,   279.1,   279.1,
  279.25,    279.25,  279.25,  279.25,
  279.5,     279.5,   279.5,   279.5,
  279.8,     279.8,   279.8,   279.8,
  280.1,     280.1,   280.1,   280.1,
  280.5,     280.5,   280.5,   280.5,
  281.05,    281.05,  281.05,  281.05,
  281.65,    281.65,  281.65,  281.65,
  282.1,     282.1,   282.1,   282.1,
  282.4,     282.4,   282.4,   282.4,
  282.65,    282.65,  282.65,  282.65,
  282.95,    282.95,  282.95,  282.95,
  283.25,    283.25,  283.25,  283.25,
  283.45,    283.45,  283.45,  283.45,
  283.55,    283.55,  283.55,  283.55,
  283.6,     283.6,   283.6,   283.6,
  283.75,    283.75,  283.75,  283.75,
  283.9,     283.9,   283.9,   283.9,
  284,       284,     284,     284,
  284.15,    284.15,  284.15,  284.15,
  284.3,     284.3,   284.3,   284.3,
  284.35,    284.35,  284.35,  284.35,
  284.4,     284.4,   284.4,   284.4,
  284.5,     284.5,   284.5,   284.5,
  284.6,     284.6,   284.6,   284.6,
  284.65,    284.65,  284.65,  284.65,
  284.65,    284.65,  284.65,  284.65,
  284.7,     284.7,   284.7,   284.7,
  284.75,    284.75,  284.75,  284.75,
  284.8,     284.8,   284.8,   284.8,
  284.9,     284.9,   284.9,   284.9,
  284.85,    284.85,  284.85,  284.85,
  284.7,     284.7,   284.7,   284.7,
  284.55,    284.55,  284.55,  284.55,
  284.4,     284.4,   284.4,   284.4,
  284.25,    284.25,  284.25,  284.25,
  284.05,    284.05,  284.05,  284.05,
  283.95,    283.95,  283.95,  283.95,
  284.1,     284.1,   284.1,   284.1,
  284.35,    284.35,  284.35,  284.35,
  284.5,     284.5,   284.5,   284.5,
  284.75,    284.75,  284.75,  284.75,
  284.95,    284.95,  284.95,  284.95,
  284.7,     284.7,   284.7,   284.7,
  284.5,     284.5,   284.5,   284.5,
  284.45,    284.45,  284.45,  284.45,
  284.15,    284.15,  284.15,  284.15,
  283.8,     283.8,   283.8,   283.8,
  283.6,     283.6,   283.6,   283.6,
  283.45,    283.45,  283.45,  283.45,
  283.2,     283.2,   283.2,   283.2,
  283,       283,     283,     283,
  282.75,    282.75,  282.75,  282.75,
  282.5,     282.5,   282.5,   282.5,
  282.4,     282.4,   282.4,   282.4,
  282.35,    282.35,  282.35,  282.35,
  282.3,     282.3,   282.3,   282.3,
  282.1,     282.1,   282.1,   282.1,
  282,       282,     282,     282,
  282.05,    282.05,  282.05,  282.05,
  282,       282,     282,     282,
  281.9,     281.9,   281.9,   281.9,
  281.9,     281.9,   281.9,   281.9,
  282,       282,     282,     282,
  282.15,    282.15,  282.15,  282.15,
  282.25,    282.25,  282.25,  282.25,
  282.3,     282.3,   282.3,   282.3,
  282.45,    282.45,  282.45,  282.45,
  282.65,    282.65,  282.65,  282.65,
  282.8,     282.8,   282.8,   282.8,
  282.95,    282.95,  282.95,  282.95,
  283.3,     283.3,   283.3,   283.3,
  283.55,    283.55,  283.55,  283.55,
  284,       284,     284,     284,
  284.6,     284.6,   284.6,   284.6,
  284.9,     284.9,   284.9,   284.9,
  285.15,    285.15,  285.15,  285.15,
  284.8,     284.8,   284.8,   284.8,
  284,       284,     284,     284,
  283.8,     283.8,   283.8,   283.8,
  283.8,     283.8,   283.8,   283.8,
  283.65,    283.65,  283.65,  283.65,
  283.6,     283.6,   283.6,   283.6,
  283.5,     283.5,   283.5,   283.5,
  283.4,     283.4,   283.4,   283.4,
  283.45,    283.45,  283.45,  283.45,
  283.6,     283.6,   283.6,   283.6,
  283.55,    283.55,  283.55,  283.55,
  283.45,    283.45,  283.45,  283.45,
  283.35,    283.35,  283.35,  283.35,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  283.15,    283.15,  283.15,  283.15,
  282.95,    282.95,  282.95,  282.95,
  282.85,    282.85,  282.85,  282.85,
  282.95,    282.95,  282.95,  282.95,
  283,       283,     283,     283,
  282.95,    282.95,  282.95,  282.95,
  282.85,    282.85,  282.85,  282.85,
  282.7,     282.7,   282.7,   282.7,
  282.7,     282.7,   282.7,   282.7,
  282.6,     282.6,   282.6,   282.6,
  282.35,    282.35,  282.35,  282.35,
  282.3,     282.3,   282.3,   282.3,
  282.1,     282.1,   282.1,   282.1,
  281.95,    281.95,  281.95,  281.95,
  281.85,    281.85,  281.85,  281.85,
  281.5,     281.5,   281.5,   281.5,
  281.25,    281.25,  281.25,  281.25,
  281.35,    281.35,  281.35,  281.35,
  281.55,    281.55,  281.55,  281.55,
  281.25,    281.25,  281.25,  281.25,
  280.85,    280.85,  280.85,  280.85,
  280.7,     280.7,   280.7,   280.7,
  280.7,     280.7,   280.7,   280.7,
  280.95,    280.95,  280.95,  280.95,
  281.15,    281.15,  281.15,  281.15,
  280.75,    280.75,  280.75,  280.75,
  280.3,     280.3,   280.3,   280.3,
  280.15,    280.15,  280.15,  280.15,
  280.05,    280.05,  280.05,  280.05,
  280.05,    280.05,  280.05,  280.05,
  279.95,    279.95,  279.95,  279.95,
  279.75,    279.75,  279.75,  279.75,
  279.5,     279.5,   279.5,   279.5,
  279.25,    279.25,  279.25,  279.25,
  279.15,    279.15,  279.15,  279.15,
  279.2,     279.2,   279.2,   279.2,
  279.25,    279.25,  279.25,  279.25,
  279.2,     279.2,   279.2,   279.2,
  279.1,     279.1,   279.1,   279.1,
  279,       279,     279,     279,
  279,       279,     279,     279,
  279.05,    279.05,  279.05,  279.05,
  278.75,    278.75,  278.75,  278.75,
  278.4,     278.4,   278.4,   278.4,
  278.3,     278.3,   278.3,   278.3,
  278.3,     278.3,   278.3,   278.3,
  278.3,     278.3,   278.3,   278.3,
  278.15,    278.15,  278.15,  278.15,
  278.1,     278.1,   278.1,   278.1,
  278.3,     278.3,   278.3,   278.3,
  278.5,     278.5,   278.5,   278.5,
  278.45,    278.45,  278.45,  278.45,
  278.15,    278.15,  278.15,  278.15,
  277.95,    277.95,  277.95,  277.95,
  278,       278,     278,     278,
  278.1,     278.1,   278.1,   278.1,
  278.25,    278.25,  278.25,  278.25,
  278.35,    278.35,  278.35,  278.35,
  278.15,    278.15,  278.15,  278.15,
  277.85,    277.85,  277.85,  277.85,
  277.85,    277.85,  277.85,  277.85,
  277.9,     277.9,   277.9,   277.9,
  277.8,     277.8,   277.8,   277.8,
  277.65,    277.65,  277.65,  277.65,
  277.45,    277.45,  277.45,  277.45,
  277.4,     277.4,   277.4,   277.4,
  277.65,    277.65,  277.65,  277.65,
  278.1,     278.1,   278.1,   278.1,
  278.55,    278.55,  278.55,  278.55,
  278.8,     278.8,   278.8,   278.8,
  278.8,     278.8,   278.8,   278.8,
  278.8,     278.8,   278.8,   278.8,
  279,       279,     279,     279,
  279.3,     279.3,   279.3,   279.3,
  279.4,     279.4,   279.4,   279.4,
  279.25,    279.25,  279.25,  279.25,
  279.2,     279.2,   279.2,   279.2,
  279.3,     279.3,   279.3,   279.3,
  279.25,    279.25,  279.25,  279.25,
  279.05,    279.05,  279.05,  279.05,
  278.95,    278.95,  278.95,  278.95,
  279.05,    279.05,  279.05,  279.05,
  279.2,     279.2,   279.2,   279.2,
  279.3,     279.3,   279.3,   279.3,
  279.3,     279.3,   279.3,   279.3,
  279.2,     279.2,   279.2,   279.2,
  279.15,    279.15,  279.15,  279.15,
  279.1,     279.1,   279.1,   279.1,
  279.05,    279.05,  279.05,  279.05,
  279,       279,     279,     279,
  278.8,     278.8,   278.8,   278.8,
  278.55,    278.55,  278.55,  278.55,
  278.4,     278.4,   278.4,   278.4,
  278.4,     278.4,   278.4,   278.4,
  278.45,    278.45,  278.45,  278.45,
  278.45,    278.45,  278.45,  278.45,
  278.4,     278.4,   278.4,   278.4,
  278.35,    278.35,  278.35,  278.35,
  278.35,    278.35,  278.35,  278.35,
  278.25,    278.25,  278.25,  278.25,
  278.1,     278.1,   278.1,   278.1,
  277.95,    277.95,  277.95,  277.95,
  277.85,    277.85,  277.85,  277.85,
  277.65,    277.65,  277.65,  277.65,
  277.35,    277.35,  277.35,  277.35,
  277.2,     277.2,   277.2,   277.2,
  277.1,     277.1,   277.1,   277.1,
  276.85,    276.85,  276.85,  276.85,
  276.55,    276.55,  276.55,  276.55,
  276.45,    276.45,  276.45,  276.45,
  276.4,     276.4,   276.4,   276.4,
  276.2,     276.2,   276.2,   276.2,
  275.95,    275.95,  275.95,  275.95,
  275.95,    275.95,  275.95,  275.95,
  276.3,     276.3,   276.3,   276.3,
  276.75,    276.75,  276.75,  276.75,
  277,       277,     277,     277,
  277.2,     277.2,   277.2,   277.2,
  277.6,     277.6,   277.6,   277.6,
  278.05,    278.05,  278.05,  278.05,
  278.45,    278.45,  278.45,  278.45,
  278.7,     278.7,   278.7,   278.7,
  278.8,     278.8,   278.8,   278.8,
  278.95,    278.95,  278.95,  278.95,
  279,       279,     279,     279,
  278.95,    278.95,  278.95,  278.95,
  278.9,     278.9,   278.9,   278.9,
  278.8,     278.8,   278.8,   278.8,
  278.65,    278.65,  278.65,  278.65,
  278.5,     278.5,   278.5,   278.5,
  278.3,     278.3,   278.3,   278.3,
  278.05,    278.05,  278.05,  278.05,
  277.9,     277.9,   277.9,   277.9,
  277.75,    277.75,  277.75,  277.75,
  277.65,    277.65,  277.65,  277.65,
  277.65,    277.65,  277.65,  277.65,
  277.6,     277.6,   277.6,   277.6,
  277.55,    277.55,  277.55,  277.55,
  277.6,     277.6,   277.6,   277.6,
  277.75,    277.75,  277.75,  277.75,
  278,       278,     278,     278,
  278.25,    278.25,  278.25,  278.25,
  278.4,     278.4,   278.4,   278.4,
  278.4,     278.4,   278.4,   278.4,
  278.25,    278.25,  278.25,  278.25,
  278.1,     278.1,   278.1,   278.1,
  278,       278,     278,     278,
  277.95,    277.95,  277.95,  277.95,
  277.9,     277.9,   277.9,   277.9,
  277.8,     277.8,   277.8,   277.8,
  277.7,     277.7,   277.7,   277.7,
  277.55,    277.55,  277.55,  277.55,
  277.5,     277.5,   277.5,   277.5,
  277.55,    277.55,  277.55,  277.55,
  277.5,     277.5,   277.5,   277.5,
  277.45,    277.45,  277.45,  277.45,
  277.2,     277.2,   277.2,   277.2,
  276.7,     276.7,   276.7,   276.7,
  276.25,    276.25,  276.25,  276.25,
  275.85,    275.85,  275.85,  275.85,
  275.65,    275.65,  275.65,  275.65,
  275.85,    275.85,  275.85,  275.85,
  276.45,    276.45,  276.45,  276.45,
  277.05,    277.05,  277.05,  277.05,
  277.55,    277.55,  277.55,  277.55,
  278.2,     278.2,   278.2,   278.2,
  278.85,    278.85,  278.85,  278.85,
  279.35,    279.35,  279.35,  279.35,
  279.6,     279.6,   279.6,   279.6,
  279.65,    279.65,  279.65,  279.65,
  279.45,    279.45,  279.45,  279.45,
  279.15,    279.15,  279.15,  279.15,
  278.85,    278.85,  278.85,  278.85,
  278.15,    278.15,  278.15,  278.15,
  277.6,     277.6,   277.6,   277.6,
  277.7,     277.7,   277.7,   277.7,
  278.05,    278.05,  278.05,  278.05,
  278.35,    278.35,  278.35,  278.35,
  278.45,    278.45,  278.45,  278.45,
  278.5,     278.5,   278.5,   278.5,
  278.55,    278.55,  278.55,  278.55,
  278.55,    278.55,  278.55,  278.55,
  278.45,    278.45,  278.45,  278.45,
  278.35,    278.35,  278.35,  278.35,
  278.25,    278.25,  278.25,  278.25,
  278.05,    278.05,  278.05,  278.05,
  277.9,     277.9,   277.9,   277.9,
  277.75,    277.75,  277.75,  277.75,
  277.5,     277.5,   277.5,   277.5,
  277.25,    277.25,  277.25,  277.25,
  277.15,    277.15,  277.15,  277.15,
  277.1,     277.1,   277.1,   277.1,
  276.85,    276.85,  276.85,  276.85,
  276.6,     276.6,   276.6,   276.6,
  276.5,     276.5,   276.5,   276.5,
  276.5,     276.5,   276.5,   276.5,
  276.5,     276.5,   276.5,   276.5,
  276.3,     276.3,   276.3,   276.3,
  276.05,    276.05,  276.05,  276.05,
  275.9,     275.9,   275.9,   275.9,
  275.9,     275.9,   275.9,   275.9,
  275.8,     275.8,   275.8,   275.8,
  275.5,     275.5,   275.5,   275.5,
  275.2,     275.2,   275.2,   275.2,
  274.95,    274.95,  274.95,  274.95,
  274.85,    274.85,  274.85,  274.85,
  274.9,     274.9,   274.9,   274.9,
  275,       275,     275,     275,
  275.1,     275.1,   275.1,   275.1,
  275.3,     275.3,   275.3,   275.3,
  275.7,     275.7,   275.7,   275.7,
  276.6,     276.6,   276.6,   276.6,
  277.6,     277.6,   277.6,   277.6,
  278.15,    278.15,  278.15,  278.15,
  278.5,     278.5,   278.5,   278.5,
  278.6,     278.6,   278.6,   278.6,
  278.6,     278.6,   278.6,   278.6,
  278.65,    278.65,  278.65,  278.65,
  278.8,     278.8,   278.8,   278.8,
  279.15,    279.15,  279.15,  279.15,
  279.45,    279.45,  279.45,  279.45,
  279.55,    279.55,  279.55,  279.55,
  279.55,    279.55,  279.55,  279.55,
  279.55,    279.55,  279.55,  279.55,
  279.65,    279.65,  279.65,  279.65,
  279.85,    279.85,  279.85,  279.85,
  280.05,    280.05,  280.05,  280.05,
  280.25,    280.25,  280.25,  280.25,
  280.4,     280.4,   280.4,   280.4,
  280.5,     280.5,   280.5,   280.5,
  280.65,    280.65,  280.65,  280.65,
  280.75,    280.75,  280.75,  280.75,
  280.75,    280.75,  280.75,  280.75,
  280.7,     280.7,   280.7,   280.7,
  280.7,     280.7,   280.7,   280.7,
  280.8,     280.8,   280.8,   280.8,
  280.85,    280.85,  280.85,  280.85,
  280.8,     280.8,   280.8,   280.8,
  280.75,    280.75,  280.75,  280.75,
  280.75,    280.75,  280.75,  280.75,
  280.8,     280.8,   280.8,   280.8,
  280.85,    280.85,  280.85,  280.85,
  280.9,     280.9,   280.9,   280.9,
  281.05,    281.05,  281.05,  281.05,
  281.2,     281.2,   281.2,   281.2,
  281.25,    281.25,  281.25,  281.25,
  281.3,     281.3,   281.3,   281.3,
  281.45,    281.45,  281.45,  281.45,
  281.5,     281.5,   281.5,   281.5,
  281.35,    281.35,  281.35,  281.35,
  281.35,    281.35,  281.35,  281.35,
  281.3,     281.3,   281.3,   281.3,
  281.15,    281.15,  281.15,  281.15,
  281,       281,     281,     281,
  280.85,    280.85,  280.85,  280.85,
  281,       281,     281,     281,
  281.2,     281.2,   281.2,   281.2,
  281.35,    281.35,  281.35,  281.35,
  281.55,    281.55,  281.55,  281.55,
  281.8,     281.8,   281.8,   281.8,
  282,       282,     282,     282,
  282.1,     282.1,   282.1,   282.1,
  282.2,     282.2,   282.2,   282.2,
  282.25,    282.25,  282.25,  282.25,
  282.25,    282.25,  282.25,  282.25,
  282.3,     282.3,   282.3,   282.3,
  282.45,    282.45,  282.45,  282.45,
  282.55,    282.55,  282.55,  282.55,
  282.55,    282.55,  282.55,  282.55,
  282.55,    282.55,  282.55,  282.55,
  282.45,    282.45,  282.45,  282.45,
  282.25,    282.25,  282.25,  282.25,
  282.05,    282.05,  282.05,  282.05,
  281.8,     281.8,   281.8,   281.8,
  281.45,    281.45,  281.45,  281.45,
  281.15,    281.15,  281.15,  281.15,
  280.95,    280.95,  280.95,  280.95,
  280.75,    280.75,  280.75,  280.75,
  280.55,    280.55,  280.55,  280.55,
  280.4,     280.4,   280.4,   280.4,
  280.3,     280.3,   280.3,   280.3,
  280.2,     280.2,   280.2,   280.2,
  280,       280,     280,     280,
  279.75,    279.75,  279.75,  279.75,
  279.6,     279.6,   279.6,   279.6,
  279.5,  279.5, 279.5,   279.5 ;

 Rainf =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0004389,
  0.0004389,
  0.0003278,
  0.0002167,
  0.0003278,
  0.0002167,
  0.0002167,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002167,
  0.0003278,
  0.0002167,
  0.0003278,
  0.0002167,
  0.0002167,
  0.0002167,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002167,
  0.0007667,
  0.0006556,
  0.0006556,
  0.0009833,
  0.0003278,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0003278,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0003278,
  0.0003278,
  0.0003278,
  0.0003278,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002167,
  0.0003278,
  0.00055,
  0.0003278,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0006556,
  0.0001111,
  0.0003278,
  0.0003278,
  0.0001111,
  0.00055,
  0.0008778,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0003278,
  0.0004389,
  0.0004389,
  0.0001111,
  0.0002167,
  0.0001111,
  0.0002167,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0.0007667,
  0.0009833,
  0.0007667,
  0.0009833,
  0.0006556,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0003278,
  0.0003278,
  0.0004389,
  0.0003278,
  0.0006556,
  0.0006556,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0004389,
  0.0001111,
  0.0001111,
  0,
  0.0004389,
  0.0002167,
  0.0003278,
  0.0008778,
  0.00055,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0006556,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0001111,
  0.0003278,
  0.0004389,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0003278,
  0.0004389,
  0.0003278,
  0.0004389,
  0.0004389,
  0.0004389,
  0.0007667,
  0.0006556,
  0.00055,
  0.0006556,
  0.0003278,
  0.0003278,
  0.0004389,
  0.0002167,
  0,
  0,
  0,
  0.0001111,
  0.0002167,
  0,
  0,
  0,
  0,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.00055,
  0.0004389,
  0.0006556,
  0.00055,
  0.00055,
  0,
  0.0003278,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0003278,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0004389,
  0.0001111,
  0,
  0,
  0.00055,
  0.0007667,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0001111,
  0.0002167,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0.0007667,
  0.0007667,
  0.001094,
  0.0001111,
  0.0001111,
  0.00055,
  0.0001111,
  0.0001111,
  0.0002167,
  0.0001111,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0.0004389,
  0,
  0,
  0,
  0.0006556,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0008778,
  0.0001111,
  0.0002167,
  0.00055,
  0.0003278,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0.0001111,
  0,
  0.0002167,
  0.0009833,
  0.00055,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0006556,
  0.0001111,
  0.0001111,
  0,
  0.0003278,
  0.0002167,
  0.0004389,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0009833,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0001111,
  0,
  0.0001111,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0.0002167,
  0.00055,
  0.0003278,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0003278,
  0.0003278,
  0.0001111,
  0,
  0.0002167,
  0.0002167,
  0.0004389,
  0.0001111,
  0.0002167,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0002167,
  0.0009833,
  0.0009833,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0008778,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0002167,
  0.0003278,
  0.0004389,
  0.0007667,
  0.0006556,
  0.0003278,
  0.0004389,
  0.00055,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0004389,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0003278,
  0,
  0.0004389,
  0.0002167,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002167,
  0.0001111,
  0.0002167,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0002167,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0.0002167,
  0.0002167,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0004389,
  0.00055,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.00055,
  0.0004389,
  0.0006556,
  0.0006556,
  0.00055,
  0.0006556,
  0.0006556,
  0.00055,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0.0001111,
  0.00055,
  0.0007667,
  0.0006556,
  0.00055,
  0.00055,
  0.0004389,
  0.0002167,
  0.0003278,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0002167,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0007667,
  0.0004389,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0006556,
  0.0009833,
  0.0004389,
  0.001094,
  0.001311,
  0.0003278,
  0.0002167,
  0,
  0.0002167,
  0,
  0.0001111,
  0.0002167,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0006556,
  0.0004389,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0001111,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.00055,
  0.0002167,
  0.0002167,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.003833,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0004389,
  0.00055,
  0.0003278,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0,
  0.0006556,
  0.0006556,
  0,
  0.0001111,
  0.0007667,
  0.0006556,
  0.0001111,
  0.0001111,
  0.0002167,
  0.0003278,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0.00055,
  0.0002167,
  0.0001111,
  0.0004389,
  0.0004389,
  0.0004389,
  0.0004389,
  0.0002167,
  0.0003278,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0004389,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0003278,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0004389,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0.0006556,
  0.0007667,
  0.00055,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002167,
  0,
  0,
  0.001311,
  0.0003278,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.00055,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0,
  0,
  0,
  0.0003278,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0002167,
  0.001533,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.001422,
  0.001533,
  0.0004389,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0004389,
  0.0002167,
  0.00055,
  0.001206,
  0.0003278,
  0.0002167,
  0.0006556,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0002167,
  0.0006556,
  0.00055,
  0.0003278,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.00055,
  0.0002167,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0004389,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0.0007667,
  0.0003278,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0004389,
  0.0003278,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.00055,
  0.0002167,
  0.0001111,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0002167,
  0.0004389,
  0.0004389,
  0.0003278,
  0.0002167,
  0.0002167,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0003278,
  0.0001111,
  0.0001111,
  0.002956,
  0.0008778,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.001094,
  0.0004389,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0004389,
  0.00055,
  0.0002167,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0003278,
  0.0004389,
  0.0002167,
  0,
  0,
  0,
  0.005472,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.001644,
  0.001206,
  0.0004389,
  0.0001111,
  0.0002167,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.00055,
  0.001422,
  0.001972,
  0.0006556,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0.00055,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0004389,
  0,
  0,
  0.0002167,
  0.0006556,
  0.0003278,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0.0002167,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0002167,
  0,
  0.0001111,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0006556,
  0.0001111,
  0.0001111,
  0.00055,
  0.0003278,
  0.0002167,
  0,
  0.0002167,
  0.0004389,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0006556,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.001644,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0002167,
  0,
  0.0004389,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.0003278,
  0.0009833,
  0.0004389,
  0.0002167,
  0.0003278,
  0.0006556,
  0.0002167,
  0.0001111,
  0.0002167,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0,
  0,
  0.0001111,
  0.0002167,
  0.0001111,
  0.0002167,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0003278,
  0.0003278,
  0.0001111,
  0.0002167,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0003278,
  0.0002167,
  0.0002167,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0.0008778,
  0.0004389,
  0.001206,
  0.002739,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0,
  0.001206,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002167,
  0.00055,
  0.0003278,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003278,
  0.00175,
  0.0009833,
  0.00175,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0006556,
  0.0002167,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.001328,
  0.0003333,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0003333,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003333,
  0.0001111,
  0,
  0.0002222,
  0.0002222,
  0.001767,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0004444,
  0.001878,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0004444,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003333,
  0.0003333,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003333,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003333,
  0,
  0.0003333,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0004444,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0006611,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003333,
  0,
  0.0008833,
  0,
  0,
  0.0004444,
  0.0004444,
  0,
  0.0002222,
  0,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.001217,
  0.0002222,
  0,
  0.0003333,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0002222,
  0.001328,
  0.00155,
  0.001767,
  0.0004444,
  0.0006611,
  0.001878,
  0.0021,
  0.0003333,
  0.0001111,
  0.001767,
  0.0007722,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0.0004444,
  0.0007722,
  0.0001111,
  0,
  0.0004444,
  0.0005556,
  0.0002222,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0004444,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0004444,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.001878,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0005556,
  0.0004444,
  0.0004444,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0002222,
  0.0002222,
  0.0003333,
  0.0003333,
  0.0003333,
  0.0001111,
  0.0001111,
  0.0002222,
  0.0004444,
  0.001217,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0003333,
  0.0001111,
  0.0001111,
  0.0004444,
  0.0001111,
  0.0001111,
  0.0002222,
  0.0003333,
  0.0002222,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0004444,
  0.0008833,
  0.001328,
  0.0003333,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0003333,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0007722,
  0.01039,
  0.001217,
  0.0004444,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.005417,
  0.0008833,
  0.001328,
  0.0021,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0002222,
  0.0002222,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0001111,
  0.0002222,
  0.001106,
  0.0009944,
  0.0005556,
  0.0007722,
  0.0008833,
  0.0007722,
  0.0007722,
  0.001106,
  0.0003333,
  0.001328,
  0.0005556,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0008833,
  0.0006611,
  0.0008833,
  0.0007722,
  0.0006611,
  0.0002222,
  0.0002222,
  0.0002222,
  0.0001111,
  0,
  0.0002222,
  0.0009944,
  0.0002222,
  0.0002222,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0005556,
  0.0003333,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.001217,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0002222,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.00155,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0004444,
  0.0007722,
  0.0006611,
  0.0004444,
  0.0003333,
  0.0003333,
  0.0003333,
  0.0003333,
  0.0006611,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0002222,
  0.0001111,
  0.0001111,
  0.0003333,
  0.0006611,
  0.0005556,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0021,
  0.0003333,
  0.0003333,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.001878,
  0,
  0,
  0,
  0.0007722,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0002222,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0003333,
  0,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0003333,
  0,
  0.0001111,
  0.0006611,
  0.0007722,
  0.0003333,
  0.0005556,
  0.0001111,
  0.0002222,
  0.0001111,
  0.0001111,
  0.0002222,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0006611,
  0.0002222,
  0,
  0.0006611,
  0.0002222,
  0.0008833,
  0.0001111,
  0.0002222,
  0.0003333,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0004444,
  0.0003333,
  0.001106,
  0.0006611,
  0.001106,
  0.0006611,
  0.0001111,
  0.0002222,
  0.0009944,
  0.003317,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0003333,
  0,
  0.0002222,
  0,
  0.0001111,
  0.0001111,
  0.0003333,
  0.0003333,
  0.0006611,
  0.0003333,
  0.0002222,
  0.0008833,
  0.0007722,
  0.0006611,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0003333,
  0.0002222,
  0,
  0.001661,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0007722,
  0.0005556,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0006611,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0.0003333,
  0.001217,
  0.0001111,
  0,
  0.0002222,
  0.0001111,
  0,
  0.0001111,
  0.0006611,
  0,
  0.0002222,
  0,
  0.0001111,
  0.0001111,
  0.0005556,
  0.0008833,
  0.0002222,
  0,
  0.0001111,
  0.0003333,
  0,
  0.0003333,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0.0002222,
  0.0005556,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0.0002222,
  0.0001111,
  0.0002222,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0004444,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0001111,
  0,
  0.0003333,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.001106,
  0.0003333,
  0.0002222,
  0.0001111,
  0.0001111,
  0,
  0.0004444,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0002222,
  0.0002222,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0005556,
  0.0003333,
  0.0004444,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003333,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0003333,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0001111,
  0.0002222,
  0.0001111,
  0.0003333,
  0.0003333,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0002222,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0003333,
  0.0002222,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0004444,
  0.0004444,
  0.0004444,
  0.0002222,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0001111,
  0.0001111,
  0.0002222,
  0.0002222,
  0.0002222,
  0.0002222,
  0.0003333,
  0.0001111,
  0.0002222,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0.0003333,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0002222,
  0.0003333,
  0.0001111,
  0.0004444,
  0.0004444,
  0.0003333,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0.0002222,
  0.0002222,
  0.0004444,
  0.0002222,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0005556,
  0.0004444,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0003333,
  0.0005556,
  0.001217,
  0.001439,
  0.0008833,
  0.0004444,
  0.0004444,
  0.0003333,
  0.0003333,
  0.0002222,
  0.0002222,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0002222,
  0.0004444,
  0.0007722,
  0.0008833,
  0.0005556,
  0.0003333,
  0.0006611,
  0.0007722,
  0.0002222,
  0.0003333,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003333,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0.0002222,
  0.0006611,
  0.0003333,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0.0002222,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0.0002222,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0002222,
  0,
  0.0001111,
  0,
  0.0002222,
  0.0006611,
  0.0002222,
  0,
  0,
  0.0002222,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0.0004444,
  0.0004444,
  0.0003333,
  0.0004444,
  0.0002222,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0004444,
  0.0001111,
  0,
  0,
  0.0002222,
  0.002767,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0.0003333,
  0.0001111,
  0,
  0,
  0.0003333,
  0.0004444,
  0.0003333,
  0,
  0,
  0,
  0.0003333,
  0.0003333,
  0.0007722,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0004444,
  0.0007722,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0003333,
  0.0001111,
  0,
  0.0006611,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0.0002222,
  0.0001111,
  0.0004444,
  0.0003333,
  0.0002222,
  0.0003333,
  0.0003333,
  0,
  0.0002222,
  0.0003333,
  0.0001111,
  0,
  0,
  0,
  0,
  0.0003333,
  0,
  0,
  0,
  0,
  0,
  0.0002222,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0.0001111,
  0.0004444,
  0.0003333,
  0.0001111,
  0.0001111,
  0,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0001111,
  0.0002222,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 Snowf =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 Qair =
  0.001384,   0.001384,    0.001384,    0.001384, 
  0.001384,   0.001384,    0.001384,    0.001384,
  0.001373,   0.001373,    0.001373,    0.001373,
  0.001362,   0.001362,    0.001362,    0.001362,
  0.001352,   0.001352,    0.001352,    0.001352,
  0.001346,   0.001346,    0.001346,    0.001346,
  0.001341,   0.001341,    0.001341,    0.001341,
  0.001335,   0.001335,    0.001335,    0.001335,
  0.001325,   0.001325,    0.001325,    0.001325,
  0.001304,   0.001304,    0.001304,    0.001304,
  0.001288,   0.001288,    0.001288,    0.001288,
  0.001283,   0.001283,    0.001283,    0.001283,
  0.001283,   0.001283,    0.001283,    0.001283,
  0.001293,   0.001293,    0.001293,    0.001293,
  0.00133,    0.00133,     0.00133,     0.00133,
  0.001361,   0.001361,    0.001361,    0.001361,
  0.001372,   0.001372,    0.001372,    0.001372,
  0.001351,   0.001351,    0.001351,    0.001351,
  0.00133,    0.00133,     0.00133,     0.00133,
  0.001357,   0.001357,    0.001357,    0.001357,
  0.001369,   0.001369,    0.001369,    0.001369,
  0.001389,   0.001389,    0.001389,    0.001389,
  0.001421,   0.001421,    0.001421,    0.001421,
  0.001431,   0.001431,    0.001431,    0.001431,
  0.001449,   0.001449,    0.001449,    0.001449,
  0.001488,   0.001488,    0.001488,    0.001488,
  0.001517,   0.001517,    0.001517,    0.001517,
  0.001533,   0.001533,    0.001533,    0.001533,
  0.001554,   0.001554,    0.001554,    0.001554,
  0.001547,   0.001547,    0.001547,    0.001547,
  0.001533,   0.001533,    0.001533,    0.001533,
  0.001558,   0.001558,    0.001558,    0.001558,
  0.00158,    0.00158,     0.00158,     0.00158,
  0.001564,   0.001564,    0.001564,    0.001564,
  0.001543,   0.001543,    0.001543,    0.001543,
  0.001501,   0.001501,    0.001501,    0.001501,
  0.001458,   0.001458,    0.001458,    0.001458,
  0.001452,   0.001452,    0.001452,    0.001452,
  0.001441,   0.001441,    0.001441,    0.001441,
  0.001412,   0.001412,    0.001412,    0.001412,
  0.001409,   0.001409,    0.001409,    0.001409,
  0.001401,   0.001401,    0.001401,    0.001401,
  0.001378,   0.001378,    0.001378,    0.001378,
  0.001361,   0.001361,    0.001361,    0.001361,
  0.001341,   0.001341,    0.001341,    0.001341,
  0.00132,    0.00132,     0.00132,     0.00132,
  0.00129,    0.00129,     0.00129,     0.00129,
  0.001275,   0.001275,    0.001275,    0.001275,
  0.00125,    0.00125,     0.00125,     0.00125,
  0.001221,   0.001221,    0.001221,    0.001221,
  0.001212,   0.001212,    0.001212,    0.001212,
  0.001207,   0.001207,    0.001207,    0.001207,
  0.001202,   0.001202,    0.001202,    0.001202,
  0.001193,   0.001193,    0.001193,    0.001193,
  0.001174,   0.001174,    0.001174,    0.001174,
  0.001151,   0.001151,    0.001151,    0.001151,
  0.001128,   0.001128,    0.001128,    0.001128,
  0.001119,   0.001119,    0.001119,    0.001119,
  0.001106,   0.001106,    0.001106,    0.001106,
  0.00108,    0.00108,     0.00108,     0.00108,
  0.001075,   0.001075,    0.001075,    0.001075,
  0.001075,   0.001075,    0.001075,    0.001075,
  0.001071,   0.001071,    0.001071,    0.001071,
  0.001071,   0.001071,    0.001071,    0.001071,
  0.001067,   0.001067,    0.001067,    0.001067,
  0.001067,   0.001067,    0.001067,    0.001067,
  0.001071,   0.001071,    0.001071,    0.001071,
  0.001106,   0.001106,    0.001106,    0.001106,
  0.001174,   0.001174,    0.001174,    0.001174,
  0.001271,   0.001271,    0.001271,    0.001271,
  0.001363,   0.001363,    0.001363,    0.001363,
  0.001435,   0.001435,    0.001435,    0.001435,
  0.001496,   0.001496,    0.001496,    0.001496,
  0.001537,   0.001537,    0.001537,    0.001537,
  0.001583,   0.001583,    0.001583,    0.001583,
  0.001594,   0.001594,    0.001594,    0.001594,
  0.001572,   0.001572,    0.001572,    0.001572,
  0.001554,   0.001554,    0.001554,    0.001554,
  0.001547,   0.001547,    0.001547,    0.001547,
  0.001551,   0.001551,    0.001551,    0.001551,
  0.001547,   0.001547,    0.001547,    0.001547,
  0.001525,   0.001525,    0.001525,    0.001525,
  0.001512,   0.001512,    0.001512,    0.001512,
  0.00152,    0.00152,     0.00152,     0.00152,
  0.001504,   0.001504,    0.001504,    0.001504,
  0.001469,   0.001469,    0.001469,    0.001469,
  0.001452,   0.001452,    0.001452,    0.001452,
  0.00144,    0.00144,     0.00144,     0.00144,
  0.001429,   0.001429,    0.001429,    0.001429,
  0.001455,   0.001455,    0.001455,    0.001455,
  0.001486,   0.001486,    0.001486,    0.001486,
  0.001486,   0.001486,    0.001486,    0.001486,
  0.001481,   0.001481,    0.001481,    0.001481,
  0.001469,   0.001469,    0.001469,    0.001469,
  0.001464,   0.001464,    0.001464,    0.001464,
  0.001469,   0.001469,    0.001469,    0.001469,
  0.001486,   0.001486,    0.001486,    0.001486,
  0.001503,   0.001503,    0.001503,    0.001503,
  0.001532,   0.001532,    0.001532,    0.001532,
  0.001585,   0.001585,    0.001585,    0.001585,
  0.001626,   0.001626,    0.001626,    0.001626,
  0.001626,   0.001626,    0.001626,    0.001626,
  0.001583,   0.001583,    0.001583,    0.001583,
  0.001545,   0.001545,    0.001545,    0.001545,
  0.001545,   0.001545,    0.001545,    0.001545,
  0.001569,   0.001569,    0.001569,    0.001569,
  0.001594,   0.001594,    0.001594,    0.001594,
  0.001606,   0.001606,    0.001606,    0.001606,
  0.0016,     0.0016,      0.0016,      0.0016,
  0.001606,   0.001606,    0.001606,    0.001606,
  0.001594,   0.001594,    0.001594,    0.001594,
  0.001575,   0.001575,    0.001575,    0.001575,
  0.001608,   0.001608,    0.001608,    0.001608,
  0.001648,   0.001648,    0.001648,    0.001648,
  0.001664,   0.001664,    0.001664,    0.001664,
  0.001673,   0.001673,    0.001673,    0.001673,
  0.001677,   0.001677,    0.001677,    0.001677,
  0.001696,   0.001696,    0.001696,    0.001696,
  0.001754,   0.001754,    0.001754,    0.001754,
  0.001822,   0.001822,    0.001822,    0.001822,
  0.001859,   0.001859,    0.001859,    0.001859,
  0.001875,   0.001875,    0.001875,    0.001875,
  0.001875,   0.001875,    0.001875,    0.001875,
  0.001876,   0.001876,    0.001876,    0.001876,
  0.001909,   0.001909,    0.001909,    0.001909,
  0.001942,   0.001942,    0.001942,    0.001942,
  0.00195,    0.00195,     0.00195,     0.00195,
  0.00195,    0.00195,     0.00195,     0.00195,
  0.001967,   0.001967,    0.001967,    0.001967,
  0.001976,   0.001976,    0.001976,    0.001976,
  0.001967,   0.001967,    0.001967,    0.001967,
  0.001959,   0.001959,    0.001959,    0.001959,
  0.001942,   0.001942,    0.001942,    0.001942,
  0.001965,   0.001965,    0.001965,    0.001965,
  0.002013,   0.002013,    0.002013,    0.002013,
  0.002039,   0.002039,    0.002039,    0.002039,
  0.002087,   0.002087,    0.002087,    0.002087,
  0.002119,   0.002119,    0.002119,    0.002119,
  0.00215,    0.00215,     0.00215,     0.00215,
  0.00219,    0.00219,     0.00219,     0.00219,
  0.002216,   0.002216,    0.002216,    0.002216,
  0.00225,    0.00225,     0.00225,     0.00225,
  0.002276,   0.002276,    0.002276,    0.002276,
  0.002285,   0.002285,    0.002285,    0.002285,
  0.002325,   0.002325,    0.002325,    0.002325,
  0.002366,   0.002366,    0.002366,    0.002366,
  0.002397,   0.002397,    0.002397,    0.002397,
  0.002429,   0.002429,    0.002429,    0.002429,
  0.002438,   0.002438,    0.002438,    0.002438,
  0.002455,   0.002455,    0.002455,    0.002455,
  0.002464,   0.002464,    0.002464,    0.002464,
  0.002464,   0.002464,    0.002464,    0.002464,
  0.002496,   0.002496,    0.002496,    0.002496,
  0.002527,   0.002527,    0.002527,    0.002527,
  0.002527,   0.002527,    0.002527,    0.002527,
  0.002496,   0.002496,    0.002496,    0.002496,
  0.002464,   0.002464,    0.002464,    0.002464,
  0.002446,   0.002446,    0.002446,    0.002446,
  0.002429,   0.002429,    0.002429,    0.002429,
  0.00242,    0.00242,     0.00242,     0.00242,
  0.002402,   0.002402,    0.002402,    0.002402,
  0.002402,   0.002402,    0.002402,    0.002402,
  0.002402,   0.002402,    0.002402,    0.002402,
  0.002385,   0.002385,    0.002385,    0.002385,
  0.002336,   0.002336,    0.002336,    0.002336,
  0.002305,   0.002305,    0.002305,    0.002305,
  0.00229,    0.00229,     0.00229,     0.00229,
  0.002268,   0.002268,    0.002268,    0.002268,
  0.002285,   0.002285,    0.002285,    0.002285,
  0.002289,   0.002289,    0.002289,    0.002289,
  0.002293,   0.002293,    0.002293,    0.002293,
  0.00232,    0.00232,     0.00232,     0.00232,
  0.002348,   0.002348,    0.002348,    0.002348,
  0.002366,   0.002366,    0.002366,    0.002366,
  0.002344,   0.002344,    0.002344,    0.002344,
  0.002321,   0.002321,    0.002321,    0.002321,
  0.002321,   0.002321,    0.002321,    0.002321,
  0.002331,   0.002331,    0.002331,    0.002331,
  0.00234,    0.00234,     0.00234,     0.00234,
  0.002349,   0.002349,    0.002349,    0.002349,
  0.002377,   0.002377,    0.002377,    0.002377,
  0.002384,   0.002384,    0.002384,    0.002384,
  0.002359,   0.002359,    0.002359,    0.002359,
  0.002357,   0.002357,    0.002357,    0.002357,
  0.002376,   0.002376,    0.002376,    0.002376,
  0.002386,   0.002386,    0.002386,    0.002386,
  0.002354,   0.002354,    0.002354,    0.002354,
  0.002294,   0.002294,    0.002294,    0.002294,
  0.002277,   0.002277,    0.002277,    0.002277,
  0.002289,   0.002289,    0.002289,    0.002289,
  0.002289,   0.002289,    0.002289,    0.002289,
  0.002248,   0.002248,    0.002248,    0.002248,
  0.002166,   0.002166,    0.002166,    0.002166,
  0.002097,   0.002097,    0.002097,    0.002097,
  0.002079,   0.002079,    0.002079,    0.002079,
  0.002097,   0.002097,    0.002097,    0.002097,
  0.002107,   0.002107,    0.002107,    0.002107,
  0.002088,   0.002088,    0.002088,    0.002088,
  0.00206,    0.00206,     0.00206,     0.00206,
  0.002082,   0.002082,    0.002082,    0.002082,
  0.002127,   0.002127,    0.002127,    0.002127,
  0.002113,   0.002113,    0.002113,    0.002113,
  0.002114,   0.002114,    0.002114,    0.002114,
  0.002179,   0.002179,    0.002179,    0.002179,
  0.002264,   0.002264,    0.002264,    0.002264,
  0.002305,   0.002305,    0.002305,    0.002305,
  0.002345,   0.002345,    0.002345,    0.002345,
  0.002402,   0.002402,    0.002402,    0.002402,
  0.00242,    0.00242,     0.00242,     0.00242,
  0.002429,   0.002429,    0.002429,    0.002429,
  0.002429,   0.002429,    0.002429,    0.002429,
  0.002406,   0.002406,    0.002406,    0.002406,
  0.00237,    0.00237,     0.00237,     0.00237,
  0.002393,   0.002393,    0.002393,    0.002393,
  0.002466,   0.002466,    0.002466,    0.002466,
  0.002481,   0.002481,    0.002481,    0.002481,
  0.00244,    0.00244,     0.00244,     0.00244,
  0.002394,   0.002394,    0.002394,    0.002394,
  0.002394,   0.002394,    0.002394,    0.002394,
  0.00245,    0.00245,     0.00245,     0.00245,
  0.002459,   0.002459,    0.002459,    0.002459,
  0.002469,   0.002469,    0.002469,    0.002469,
  0.002485,   0.002485,    0.002485,    0.002485,
  0.002473,   0.002473,    0.002473,    0.002473,
  0.002507,   0.002507,    0.002507,    0.002507,
  0.002498,   0.002498,    0.002498,    0.002498,
  0.002447,   0.002447,    0.002447,    0.002447,
  0.002436,   0.002436,    0.002436,    0.002436,
  0.0024,     0.0024,      0.0024,      0.0024,
  0.002318,   0.002318,    0.002318,    0.002318,
  0.002253,   0.002253,    0.002253,    0.002253,
  0.0022,     0.0022,      0.0022,      0.0022,
  0.002125,   0.002125,    0.002125,    0.002125,
  0.002081,   0.002081,    0.002081,    0.002081,
  0.002073,   0.002073,    0.002073,    0.002073,
  0.002045,   0.002045,    0.002045,    0.002045,
  0.001995,   0.001995,    0.001995,    0.001995,
  0.001947,   0.001947,    0.001947,    0.001947,
  0.001947,   0.001947,    0.001947,    0.001947,
  0.001988,   0.001988,    0.001988,    0.001988,
  0.002009,   0.002009,    0.002009,    0.002009,
  0.001995,   0.001995,    0.001995,    0.001995,
  0.001961,   0.001961,    0.001961,    0.001961,
  0.001982,   0.001982,    0.001982,    0.001982,
  0.002059,   0.002059,    0.002059,    0.002059,
  0.002147,   0.002147,    0.002147,    0.002147,
  0.002262,   0.002262,    0.002262,    0.002262,
  0.002381,   0.002381,    0.002381,    0.002381,
  0.002446,   0.002446,    0.002446,    0.002446,
  0.002463,   0.002463,    0.002463,    0.002463,
  0.002446,   0.002446,    0.002446,    0.002446,
  0.00243,    0.00243,     0.00243,     0.00243,
  0.002413,   0.002413,    0.002413,    0.002413,
  0.00238,    0.00238,     0.00238,     0.00238,
  0.002356,   0.002356,    0.002356,    0.002356,
  0.00234,    0.00234,     0.00234,     0.00234,
  0.002332,   0.002332,    0.002332,    0.002332,
  0.00234,    0.00234,     0.00234,     0.00234,
  0.002332,   0.002332,    0.002332,    0.002332,
  0.002245,   0.002245,    0.002245,    0.002245,
  0.002167,   0.002167,    0.002167,    0.002167,
  0.002144,   0.002144,    0.002144,    0.002144,
  0.002121,   0.002121,    0.002121,    0.002121,
  0.002129,   0.002129,    0.002129,    0.002129,
  0.002128,   0.002128,    0.002128,    0.002128,
  0.002065,   0.002065,    0.002065,    0.002065,
  0.00197,    0.00197,     0.00197,     0.00197,
  0.001899,   0.001899,    0.001899,    0.001899,
  0.001875,   0.001875,    0.001875,    0.001875,
  0.001914,   0.001914,    0.001914,    0.001914,
  0.001938,   0.001938,    0.001938,    0.001938,
  0.001907,   0.001907,    0.001907,    0.001907,
  0.001908,   0.001908,    0.001908,    0.001908,
  0.001934,   0.001934,    0.001934,    0.001934,
  0.001952,   0.001952,    0.001952,    0.001952,
  0.001993,   0.001993,    0.001993,    0.001993,
  0.002025,   0.002025,    0.002025,    0.002025,
  0.002025,   0.002025,    0.002025,    0.002025,
  0.002049,   0.002049,    0.002049,    0.002049,
  0.002059,   0.002059,    0.002059,    0.002059,
  0.002038,   0.002038,    0.002038,    0.002038,
  0.002045,   0.002045,    0.002045,    0.002045,
  0.002103,   0.002103,    0.002103,    0.002103,
  0.002185,   0.002185,    0.002185,    0.002185,
  0.002253,   0.002253,    0.002253,    0.002253,
  0.002316,   0.002316,    0.002316,    0.002316,
  0.002356,   0.002356,    0.002356,    0.002356,
  0.00238,    0.00238,     0.00238,     0.00238,
  0.002405,   0.002405,    0.002405,    0.002405,
  0.00239,    0.00239,     0.00239,     0.00239,
  0.002367,   0.002367,    0.002367,    0.002367,
  0.002375,   0.002375,    0.002375,    0.002375,
  0.002391,   0.002391,    0.002391,    0.002391,
  0.002417,   0.002417,    0.002417,    0.002417,
  0.002419,   0.002419,    0.002419,    0.002419,
  0.002422,   0.002422,    0.002422,    0.002422,
  0.002448,   0.002448,    0.002448,    0.002448,
  0.002443,   0.002443,    0.002443,    0.002443,
  0.002438,   0.002438,    0.002438,    0.002438,
  0.002455,   0.002455,    0.002455,    0.002455,
  0.002473,   0.002473,    0.002473,    0.002473,
  0.002491,   0.002491,    0.002491,    0.002491,
  0.002518,   0.002518,    0.002518,    0.002518,
  0.002546,   0.002546,    0.002546,    0.002546,
  0.002514,   0.002514,    0.002514,    0.002514,
  0.002455,   0.002455,    0.002455,    0.002455,
  0.002437,   0.002437,    0.002437,    0.002437,
  0.002446,   0.002446,    0.002446,    0.002446,
  0.002464,   0.002464,    0.002464,    0.002464,
  0.002492,   0.002492,    0.002492,    0.002492,
  0.002488,   0.002488,    0.002488,    0.002488,
  0.002475,   0.002475,    0.002475,    0.002475,
  0.002485,   0.002485,    0.002485,    0.002485,
  0.002485,   0.002485,    0.002485,    0.002485,
  0.002453,   0.002453,    0.002453,    0.002453,
  0.00244,    0.00244,     0.00244,     0.00244,
  0.002447,   0.002447,    0.002447,    0.002447,
  0.002444,   0.002444,    0.002444,    0.002444,
  0.002444,   0.002444,    0.002444,    0.002444,
  0.002466,   0.002466,    0.002466,    0.002466,
  0.002469,   0.002469,    0.002469,    0.002469,
  0.002466,   0.002466,    0.002466,    0.002466,
  0.002496,   0.002496,    0.002496,    0.002496,
  0.002473,   0.002473,    0.002473,    0.002473,
  0.002452,   0.002452,    0.002452,    0.002452,
  0.002437,   0.002437,    0.002437,    0.002437,
  0.002382,   0.002382,    0.002382,    0.002382,
  0.002332,   0.002332,    0.002332,    0.002332,
  0.0023,     0.0023,      0.0023,      0.0023,
  0.002253,   0.002253,    0.002253,    0.002253,
  0.002253,   0.002253,    0.002253,    0.002253,
  0.002324,   0.002324,    0.002324,    0.002324,
  0.002389,   0.002389,    0.002389,    0.002389,
  0.002405,   0.002405,    0.002405,    0.002405,
  0.00238,    0.00238,     0.00238,     0.00238,
  0.002364,   0.002364,    0.002364,    0.002364,
  0.002364,   0.002364,    0.002364,    0.002364,
  0.002364,   0.002364,    0.002364,    0.002364,
  0.002356,   0.002356,    0.002356,    0.002356,
  0.002324,   0.002324,    0.002324,    0.002324,
  0.002284,   0.002284,    0.002284,    0.002284,
  0.002261,   0.002261,    0.002261,    0.002261,
  0.002238,   0.002238,    0.002238,    0.002238,
  0.002207,   0.002207,    0.002207,    0.002207,
  0.002184,   0.002184,    0.002184,    0.002184,
  0.002169,   0.002169,    0.002169,    0.002169,
  0.002162,   0.002162,    0.002162,    0.002162,
  0.002154,   0.002154,    0.002154,    0.002154,
  0.002132,   0.002132,    0.002132,    0.002132,
  0.00211,    0.00211,     0.00211,     0.00211,
  0.002095,   0.002095,    0.002095,    0.002095,
  0.002095,   0.002095,    0.002095,    0.002095,
  0.00211,    0.00211,     0.00211,     0.00211,
  0.002125,   0.002125,    0.002125,    0.002125,
  0.002139,   0.002139,    0.002139,    0.002139,
  0.002147,   0.002147,    0.002147,    0.002147,
  0.002154,   0.002154,    0.002154,    0.002154,
  0.002169,   0.002169,    0.002169,    0.002169,
  0.002177,   0.002177,    0.002177,    0.002177,
  0.002177,   0.002177,    0.002177,    0.002177,
  0.002184,   0.002184,    0.002184,    0.002184,
  0.002207,   0.002207,    0.002207,    0.002207,
  0.002206,   0.002206,    0.002206,    0.002206,
  0.002198,   0.002198,    0.002198,    0.002198,
  0.002206,   0.002206,    0.002206,    0.002206,
  0.002221,   0.002221,    0.002221,    0.002221,
  0.002214,   0.002214,    0.002214,    0.002214,
  0.00219,    0.00219,     0.00219,     0.00219,
  0.002198,   0.002198,    0.002198,    0.002198,
  0.002198,   0.002198,    0.002198,    0.002198,
  0.002152,   0.002152,    0.002152,    0.002152,
  0.002106,   0.002106,    0.002106,    0.002106,
  0.002075,   0.002075,    0.002075,    0.002075,
  0.002036,   0.002036,    0.002036,    0.002036,
  0.002013,   0.002013,    0.002013,    0.002013,
  0.00203,    0.00203,     0.00203,     0.00203,
  0.00204,    0.00204,     0.00204,     0.00204,
  0.002018,   0.002018,    0.002018,    0.002018,
  0.002018,   0.002018,    0.002018,    0.002018,
  0.002025,   0.002025,    0.002025,    0.002025,
  0.002025,   0.002025,    0.002025,    0.002025,
  0.002011,   0.002011,    0.002011,    0.002011,
  0.001989,   0.001989,    0.001989,    0.001989,
  0.001968,   0.001968,    0.001968,    0.001968,
  0.001953,   0.001953,    0.001953,    0.001953,
  0.001978,   0.001978,    0.001978,    0.001978,
  0.001971,   0.001971,    0.001971,    0.001971,
  0.001932,   0.001932,    0.001932,    0.001932,
  0.001957,   0.001957,    0.001957,    0.001957,
  0.001964,   0.001964,    0.001964,    0.001964,
  0.001964,   0.001964,    0.001964,    0.001964,
  0.001988,   0.001988,    0.001988,    0.001988,
  0.001957,   0.001957,    0.001957,    0.001957,
  0.00195,    0.00195,     0.00195,     0.00195,
  0.001974,   0.001974,    0.001974,    0.001974,
  0.001968,   0.001968,    0.001968,    0.001968,
  0.001954,   0.001954,    0.001954,    0.001954,
  0.00194,    0.00194,     0.00194,     0.00194,
  0.001947,   0.001947,    0.001947,    0.001947,
  0.001989,   0.001989,    0.001989,    0.001989,
  0.002045,   0.002045,    0.002045,    0.002045,
  0.002088,   0.002088,    0.002088,    0.002088,
  0.00211,    0.00211,     0.00211,     0.00211,
  0.002117,   0.002117,    0.002117,    0.002117,
  0.002125,   0.002125,    0.002125,    0.002125,
  0.002147,   0.002147,    0.002147,    0.002147,
  0.002145,   0.002145,    0.002145,    0.002145,
  0.002152,   0.002152,    0.002152,    0.002152,
  0.002159,   0.002159,    0.002159,    0.002159,
  0.002166,   0.002166,    0.002166,    0.002166,
  0.002198,   0.002198,    0.002198,    0.002198,
  0.002174,   0.002174,    0.002174,    0.002174,
  0.002159,   0.002159,    0.002159,    0.002159,
  0.002175,   0.002175,    0.002175,    0.002175,
  0.002175,   0.002175,    0.002175,    0.002175,
  0.002175,   0.002175,    0.002175,    0.002175,
  0.002167,   0.002167,    0.002167,    0.002167,
  0.002143,   0.002143,    0.002143,    0.002143,
  0.002127,   0.002127,    0.002127,    0.002127,
  0.002143,   0.002143,    0.002143,    0.002143,
  0.002191,   0.002191,    0.002191,    0.002191,
  0.002289,   0.002289,    0.002289,    0.002289,
  0.002379,   0.002379,    0.002379,    0.002379,
  0.002453,   0.002453,    0.002453,    0.002453,
  0.002511,   0.002511,    0.002511,    0.002511,
  0.002506,   0.002506,    0.002506,    0.002506,
  0.002509,   0.002509,    0.002509,    0.002509,
  0.002545,   0.002545,    0.002545,    0.002545,
  0.002591,   0.002591,    0.002591,    0.002591,
  0.002636,   0.002636,    0.002636,    0.002636,
  0.002655,   0.002655,    0.002655,    0.002655,
  0.002633,   0.002633,    0.002633,    0.002633,
  0.00262,    0.00262,     0.00262,     0.00262,
  0.002648,   0.002648,    0.002648,    0.002648,
  0.002645,   0.002645,    0.002645,    0.002645,
  0.002633,   0.002633,    0.002633,    0.002633,
  0.002674,   0.002674,    0.002674,    0.002674,
  0.002715,   0.002715,    0.002715,    0.002715,
  0.002735,   0.002735,    0.002735,    0.002735,
  0.002744,   0.002744,    0.002744,    0.002744,
  0.002735,   0.002735,    0.002735,    0.002735,
  0.002725,   0.002725,    0.002725,    0.002725,
  0.002693,   0.002693,    0.002693,    0.002693,
  0.002599,   0.002599,    0.002599,    0.002599,
  0.002536,   0.002536,    0.002536,    0.002536,
  0.002526,   0.002526,    0.002526,    0.002526,
  0.002475,   0.002475,    0.002475,    0.002475,
  0.002434,   0.002434,    0.002434,    0.002434,
  0.002434,   0.002434,    0.002434,    0.002434,
  0.002425,   0.002425,    0.002425,    0.002425,
  0.002437,   0.002437,    0.002437,    0.002437,
  0.002469,   0.002469,    0.002469,    0.002469,
  0.002469,   0.002469,    0.002469,    0.002469,
  0.002491,   0.002491,    0.002491,    0.002491,
  0.002576,   0.002576,    0.002576,    0.002576,
  0.002661,   0.002661,    0.002661,    0.002661,
  0.002724,   0.002724,    0.002724,    0.002724,
  0.002774,   0.002774,    0.002774,    0.002774,
  0.002759,   0.002759,    0.002759,    0.002759,
  0.002672,   0.002672,    0.002672,    0.002672,
  0.002543,   0.002543,    0.002543,    0.002543,
  0.002478,   0.002478,    0.002478,    0.002478,
  0.002478,   0.002478,    0.002478,    0.002478,
  0.0025,     0.0025,      0.0025,      0.0025,
  0.002532,   0.002532,    0.002532,    0.002532,
  0.002532,   0.002532,    0.002532,    0.002532,
  0.002532,   0.002532,    0.002532,    0.002532,
  0.002522,   0.002522,    0.002522,    0.002522,
  0.002522,   0.002522,    0.002522,    0.002522,
  0.002532,   0.002532,    0.002532,    0.002532,
  0.002532,   0.002532,    0.002532,    0.002532,
  0.002541,   0.002541,    0.002541,    0.002541,
  0.002541,   0.002541,    0.002541,    0.002541,
  0.002541,   0.002541,    0.002541,    0.002541,
  0.002541,   0.002541,    0.002541,    0.002541,
  0.002541,   0.002541,    0.002541,    0.002541,
  0.002541,   0.002541,    0.002541,    0.002541,
  0.002541,   0.002541,    0.002541,    0.002541,
  0.002551,   0.002551,    0.002551,    0.002551,
  0.002583,   0.002583,    0.002583,    0.002583,
  0.002604,   0.002604,    0.002604,    0.002604,
  0.002563,   0.002563,    0.002563,    0.002563,
  0.002532,   0.002532,    0.002532,    0.002532,
  0.002553,   0.002553,    0.002553,    0.002553,
  0.002565,   0.002565,    0.002565,    0.002565,
  0.002565,   0.002565,    0.002565,    0.002565,
  0.002534,   0.002534,    0.002534,    0.002534,
  0.002483,   0.002483,    0.002483,    0.002483,
  0.002463,   0.002463,    0.002463,    0.002463,
  0.002444,   0.002444,    0.002444,    0.002444,
  0.002434,   0.002434,    0.002434,    0.002434,
  0.002434,   0.002434,    0.002434,    0.002434,
  0.002425,   0.002425,    0.002425,    0.002425,
  0.002447,   0.002447,    0.002447,    0.002447,
  0.002478,   0.002478,    0.002478,    0.002478,
  0.002469,   0.002469,    0.002469,    0.002469,
  0.002469,   0.002469,    0.002469,    0.002469,
  0.002478,   0.002478,    0.002478,    0.002478,
  0.002456,   0.002456,    0.002456,    0.002456,
  0.002454,   0.002454,    0.002454,    0.002454,
  0.002492,   0.002492,    0.002492,    0.002492,
  0.002532,   0.002532,    0.002532,    0.002532,
  0.00253,    0.00253,     0.00253,     0.00253,
  0.00254,    0.00254,     0.00254,     0.00254,
  0.002571,   0.002571,    0.002571,    0.002571,
  0.002571,   0.002571,    0.002571,    0.002571,
  0.00255,    0.00255,     0.00255,     0.00255,
  0.002538,   0.002538,    0.002538,    0.002538,
  0.002538,   0.002538,    0.002538,    0.002538,
  0.002507,   0.002507,    0.002507,    0.002507,
  0.002517,   0.002517,    0.002517,    0.002517,
  0.002517,   0.002517,    0.002517,    0.002517,
  0.002455,   0.002455,    0.002455,    0.002455,
  0.002447,   0.002447,    0.002447,    0.002447,
  0.00249,    0.00249,     0.00249,     0.00249,
  0.002502,   0.002502,    0.002502,    0.002502,
  0.002514,   0.002514,    0.002514,    0.002514,
  0.002526,   0.002526,    0.002526,    0.002526,
  0.002538,   0.002538,    0.002538,    0.002538,
  0.002532,   0.002532,    0.002532,    0.002532,
  0.002488,   0.002488,    0.002488,    0.002488,
  0.0025,     0.0025,      0.0025,      0.0025,
  0.002501,   0.002501,    0.002501,    0.002501,
  0.002479,   0.002479,    0.002479,    0.002479,
  0.002459,   0.002459,    0.002459,    0.002459,
  0.002465,   0.002465,    0.002465,    0.002465,
  0.002474,   0.002474,    0.002474,    0.002474,
  0.002491,   0.002491,    0.002491,    0.002491,
  0.002508,   0.002508,    0.002508,    0.002508,
  0.002499,   0.002499,    0.002499,    0.002499,
  0.002505,   0.002505,    0.002505,    0.002505,
  0.002497,   0.002497,    0.002497,    0.002497,
  0.002497,   0.002497,    0.002497,    0.002497,
  0.002488,   0.002488,    0.002488,    0.002488,
  0.002488,   0.002488,    0.002488,    0.002488,
  0.002499,   0.002499,    0.002499,    0.002499,
  0.002546,   0.002546,    0.002546,    0.002546,
  0.002586,   0.002586,    0.002586,    0.002586,
  0.002577,   0.002577,    0.002577,    0.002577,
  0.00257,    0.00257,     0.00257,     0.00257,
  0.002585,   0.002585,    0.002585,    0.002585,
  0.002614,   0.002614,    0.002614,    0.002614,
  0.002601,   0.002601,    0.002601,    0.002601,
  0.002589,   0.002589,    0.002589,    0.002589,
  0.002618,   0.002618,    0.002618,    0.002618,
  0.002648,   0.002648,    0.002648,    0.002648,
  0.002677,   0.002677,    0.002677,    0.002677,
  0.002686,   0.002686,    0.002686,    0.002686,
  0.002715,   0.002715,    0.002715,    0.002715,
  0.002819,   0.002819,    0.002819,    0.002819,
  0.002958,   0.002958,    0.002958,    0.002958,
  0.003091,   0.003091,    0.003091,    0.003091,
  0.003253,   0.003253,    0.003253,    0.003253,
  0.003469,   0.003469,    0.003469,    0.003469,
  0.003594,   0.003594,    0.003594,    0.003594,
  0.003628,   0.003628,    0.003628,    0.003628,
  0.00367,    0.00367,     0.00367,     0.00367,
  0.003707,   0.003707,    0.003707,    0.003707,
  0.003713,   0.003713,    0.003713,    0.003713,
  0.003732,   0.003732,    0.003732,    0.003732,
  0.003802,   0.003802,    0.003802,    0.003802,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003991,   0.003991,    0.003991,    0.003991,
  0.004054,   0.004054,    0.004054,    0.004054,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004176,   0.004176,    0.004176,    0.004176,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004128,   0.004128,    0.004128,    0.004128,
  0.003656,   0.003656,    0.003656,    0.003656,
  0.003297,   0.003297,    0.003297,    0.003297,
  0.003172,   0.003172,    0.003172,    0.003172,
  0.003148,   0.003148,    0.003148,    0.003148,
  0.003177,   0.003177,    0.003177,    0.003177,
  0.00319,    0.00319,     0.00319,     0.00319,
  0.00318,    0.00318,     0.00318,     0.00318,
  0.003193,   0.003193,    0.003193,    0.003193,
  0.003229,   0.003229,    0.003229,    0.003229,
  0.003244,   0.003244,    0.003244,    0.003244,
  0.00325,    0.00325,     0.00325,     0.00325,
  0.00328,    0.00328,     0.00328,     0.00328,
  0.003313,   0.003313,    0.003313,    0.003313,
  0.003319,   0.003319,    0.003319,    0.003319,
  0.0033,     0.0033,      0.0033,      0.0033,
  0.003328,   0.003328,    0.003328,    0.003328,
  0.00338,    0.00338,     0.00338,     0.00338,
  0.003412,   0.003412,    0.003412,    0.003412,
  0.003461,   0.003461,    0.003461,    0.003461,
  0.003549,   0.003549,    0.003549,    0.003549,
  0.003661,   0.003661,    0.003661,    0.003661,
  0.00372,    0.00372,     0.00372,     0.00372,
  0.003717,   0.003717,    0.003717,    0.003717,
  0.003683,   0.003683,    0.003683,    0.003683,
  0.003644,   0.003644,    0.003644,    0.003644,
  0.003619,   0.003619,    0.003619,    0.003619,
  0.0036,     0.0036,      0.0036,      0.0036,
  0.003581,   0.003581,    0.003581,    0.003581,
  0.003556,   0.003556,    0.003556,    0.003556,
  0.003531,   0.003531,    0.003531,    0.003531,
  0.003514,   0.003514,    0.003514,    0.003514,
  0.003497,   0.003497,    0.003497,    0.003497,
  0.003485,   0.003485,    0.003485,    0.003485,
  0.003473,   0.003473,    0.003473,    0.003473,
  0.003449,   0.003449,    0.003449,    0.003449,
  0.003413,   0.003413,    0.003413,    0.003413,
  0.00337,    0.00337,     0.00337,     0.00337,
  0.003342,   0.003342,    0.003342,    0.003342,
  0.003319,   0.003319,    0.003319,    0.003319,
  0.003311,   0.003311,    0.003311,    0.003311,
  0.003308,   0.003308,    0.003308,    0.003308,
  0.003233,   0.003233,    0.003233,    0.003233,
  0.003154,   0.003154,    0.003154,    0.003154,
  0.00312,    0.00312,     0.00312,     0.00312,
  0.003031,   0.003031,    0.003031,    0.003031,
  0.002895,   0.002895,    0.002895,    0.002895,
  0.002764,   0.002764,    0.002764,    0.002764,
  0.00259,    0.00259,     0.00259,     0.00259,
  0.002475,   0.002475,    0.002475,    0.002475,
  0.002414,   0.002414,    0.002414,    0.002414,
  0.00214,    0.00214,     0.00214,     0.00214,
  0.001806,   0.001806,    0.001806,    0.001806,
  0.001712,   0.001712,    0.001712,    0.001712,
  0.001732,   0.001732,    0.001732,    0.001732,
  0.001829,   0.001829,    0.001829,    0.001829,
  0.002018,   0.002018,    0.002018,    0.002018,
  0.00212,    0.00212,     0.00212,     0.00212,
  0.002183,   0.002183,    0.002183,    0.002183,
  0.002266,   0.002266,    0.002266,    0.002266,
  0.002339,   0.002339,    0.002339,    0.002339,
  0.002366,   0.002366,    0.002366,    0.002366,
  0.002351,   0.002351,    0.002351,    0.002351,
  0.002369,   0.002369,    0.002369,    0.002369,
  0.002392,   0.002392,    0.002392,    0.002392,
  0.002452,   0.002452,    0.002452,    0.002452,
  0.002521,   0.002521,    0.002521,    0.002521,
  0.002563,   0.002563,    0.002563,    0.002563,
  0.002627,   0.002627,    0.002627,    0.002627,
  0.002681,   0.002681,    0.002681,    0.002681,
  0.002712,   0.002712,    0.002712,    0.002712,
  0.00277,    0.00277,     0.00277,     0.00277,
  0.002835,   0.002835,    0.002835,    0.002835,
  0.002891,   0.002891,    0.002891,    0.002891,
  0.00294,    0.00294,     0.00294,     0.00294,
  0.002935,   0.002935,    0.002935,    0.002935,
  0.002913,   0.002913,    0.002913,    0.002913,
  0.002917,   0.002917,    0.002917,    0.002917,
  0.002922,   0.002922,    0.002922,    0.002922,
  0.002916,   0.002916,    0.002916,    0.002916,
  0.002879,   0.002879,    0.002879,    0.002879,
  0.002866,   0.002866,    0.002866,    0.002866,
  0.002864,   0.002864,    0.002864,    0.002864,
  0.002852,   0.002852,    0.002852,    0.002852,
  0.002841,   0.002841,    0.002841,    0.002841,
  0.002787,   0.002787,    0.002787,    0.002787,
  0.002777,   0.002777,    0.002777,    0.002777,
  0.002777,   0.002777,    0.002777,    0.002777,
  0.002746,   0.002746,    0.002746,    0.002746,
  0.002747,   0.002747,    0.002747,    0.002747,
  0.002747,   0.002747,    0.002747,    0.002747,
  0.002736,   0.002736,    0.002736,    0.002736,
  0.002745,   0.002745,    0.002745,    0.002745,
  0.002768,   0.002768,    0.002768,    0.002768,
  0.002809,   0.002809,    0.002809,    0.002809,
  0.002857,   0.002857,    0.002857,    0.002857,
  0.002877,   0.002877,    0.002877,    0.002877,
  0.002892,   0.002892,    0.002892,    0.002892,
  0.002926,   0.002926,    0.002926,    0.002926,
  0.002956,   0.002956,    0.002956,    0.002956,
  0.002991,   0.002991,    0.002991,    0.002991,
  0.00303,    0.00303,     0.00303,     0.00303,
  0.003059,   0.003059,    0.003059,    0.003059,
  0.003075,   0.003075,    0.003075,    0.003075,
  0.003091,   0.003091,    0.003091,    0.003091,
  0.003091,   0.003091,    0.003091,    0.003091,
  0.003095,   0.003095,    0.003095,    0.003095,
  0.003129,   0.003129,    0.003129,    0.003129,
  0.003146,   0.003146,    0.003146,    0.003146,
  0.003149,   0.003149,    0.003149,    0.003149,
  0.003119,   0.003119,    0.003119,    0.003119,
  0.003109,   0.003109,    0.003109,    0.003109,
  0.003134,   0.003134,    0.003134,    0.003134,
  0.003143,   0.003143,    0.003143,    0.003143,
  0.003141,   0.003141,    0.003141,    0.003141,
  0.00313,    0.00313,     0.00313,     0.00313,
  0.003086,   0.003086,    0.003086,    0.003086,
  0.003074,   0.003074,    0.003074,    0.003074,
  0.003074,   0.003074,    0.003074,    0.003074,
  0.003019,   0.003019,    0.003019,    0.003019,
  0.002996,   0.002996,    0.002996,    0.002996,
  0.002984,   0.002984,    0.002984,    0.002984,
  0.002953,   0.002953,    0.002953,    0.002953,
  0.00295,    0.00295,     0.00295,     0.00295,
  0.002932,   0.002932,    0.002932,    0.002932,
  0.002905,   0.002905,    0.002905,    0.002905,
  0.002903,   0.002903,    0.002903,    0.002903,
  0.002903,   0.002903,    0.002903,    0.002903,
  0.002914,   0.002914,    0.002914,    0.002914,
  0.002924,   0.002924,    0.002924,    0.002924,
  0.002903,   0.002903,    0.002903,    0.002903,
  0.002893,   0.002893,    0.002893,    0.002893,
  0.002874,   0.002874,    0.002874,    0.002874,
  0.002865,   0.002865,    0.002865,    0.002865,
  0.002896,   0.002896,    0.002896,    0.002896,
  0.002896,   0.002896,    0.002896,    0.002896,
  0.002876,   0.002876,    0.002876,    0.002876,
  0.002847,   0.002847,    0.002847,    0.002847,
  0.002827,   0.002827,    0.002827,    0.002827,
  0.002857,   0.002857,    0.002857,    0.002857,
  0.002894,   0.002894,    0.002894,    0.002894,
  0.002947,   0.002947,    0.002947,    0.002947,
  0.003056,   0.003056,    0.003056,    0.003056,
  0.003163,   0.003163,    0.003163,    0.003163,
  0.003219,   0.003219,    0.003219,    0.003219,
  0.003281,   0.003281,    0.003281,    0.003281,
  0.003313,   0.003313,    0.003313,    0.003313,
  0.003326,   0.003326,    0.003326,    0.003326,
  0.00333,    0.00333,     0.00333,     0.00333,
  0.003319,   0.003319,    0.003319,    0.003319,
  0.003331,   0.003331,    0.003331,    0.003331,
  0.003291,   0.003291,    0.003291,    0.003291,
  0.003286,   0.003286,    0.003286,    0.003286,
  0.003329,   0.003329,    0.003329,    0.003329,
  0.003335,   0.003335,    0.003335,    0.003335,
  0.003302,   0.003302,    0.003302,    0.003302,
  0.003255,   0.003255,    0.003255,    0.003255,
  0.003235,   0.003235,    0.003235,    0.003235,
  0.003221,   0.003221,    0.003221,    0.003221,
  0.003204,   0.003204,    0.003204,    0.003204,
  0.003165,   0.003165,    0.003165,    0.003165,
  0.003146,   0.003146,    0.003146,    0.003146,
  0.003153,   0.003153,    0.003153,    0.003153,
  0.003147,   0.003147,    0.003147,    0.003147,
  0.00314,    0.00314,     0.00314,     0.00314,
  0.003153,   0.003153,    0.003153,    0.003153,
  0.003167,   0.003167,    0.003167,    0.003167,
  0.003143,   0.003143,    0.003143,    0.003143,
  0.00315,    0.00315,     0.00315,     0.00315,
  0.003158,   0.003158,    0.003158,    0.003158,
  0.003153,   0.003153,    0.003153,    0.003153,
  0.003161,   0.003161,    0.003161,    0.003161,
  0.003134,   0.003134,    0.003134,    0.003134,
  0.003107,   0.003107,    0.003107,    0.003107,
  0.003087,   0.003087,    0.003087,    0.003087,
  0.003076,   0.003076,    0.003076,    0.003076,
  0.003087,   0.003087,    0.003087,    0.003087,
  0.003067,   0.003067,    0.003067,    0.003067,
  0.003048,   0.003048,    0.003048,    0.003048,
  0.003039,   0.003039,    0.003039,    0.003039,
  0.003036,   0.003036,    0.003036,    0.003036,
  0.003056,   0.003056,    0.003056,    0.003056,
  0.003059,   0.003059,    0.003059,    0.003059,
  0.003039,   0.003039,    0.003039,    0.003039,
  0.003024,   0.003024,    0.003024,    0.003024,
  0.00301,    0.00301,     0.00301,     0.00301,
  0.00301,    0.00301,     0.00301,     0.00301,
  0.00304,    0.00304,     0.00304,     0.00304,
  0.003087,   0.003087,    0.003087,    0.003087,
  0.003122,   0.003122,    0.003122,    0.003122,
  0.003174,   0.003174,    0.003174,    0.003174,
  0.003261,   0.003261,    0.003261,    0.003261,
  0.003299,   0.003299,    0.003299,    0.003299,
  0.003302,   0.003302,    0.003302,    0.003302,
  0.003286,   0.003286,    0.003286,    0.003286,
  0.003257,   0.003257,    0.003257,    0.003257,
  0.003247,   0.003247,    0.003247,    0.003247,
  0.003249,   0.003249,    0.003249,    0.003249,
  0.00326,    0.00326,     0.00326,     0.00326,
  0.003278,   0.003278,    0.003278,    0.003278,
  0.003317,   0.003317,    0.003317,    0.003317,
  0.00336,    0.00336,     0.00336,     0.00336,
  0.00338,    0.00338,     0.00338,     0.00338,
  0.003422,   0.003422,    0.003422,    0.003422,
  0.003426,   0.003426,    0.003426,    0.003426,
  0.003406,   0.003406,    0.003406,    0.003406,
  0.003453,   0.003453,    0.003453,    0.003453,
  0.0035,     0.0035,      0.0035,      0.0035,
  0.003547,   0.003547,    0.003547,    0.003547,
  0.00361,    0.00361,     0.00361,     0.00361,
  0.003657,   0.003657,    0.003657,    0.003657,
  0.003752,   0.003752,    0.003752,    0.003752,
  0.003913,   0.003913,    0.003913,    0.003913,
  0.004043,   0.004043,    0.004043,    0.004043,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004172,   0.004172,    0.004172,    0.004172,
  0.004217,   0.004217,    0.004217,    0.004217,
  0.004278,   0.004278,    0.004278,    0.004278,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.004689,   0.004689,    0.004689,    0.004689,
  0.004956,   0.004956,    0.004956,    0.004956,
  0.005048,   0.005048,    0.005048,    0.005048,
  0.005078,   0.005078,    0.005078,    0.005078,
  0.00514,    0.00514,     0.00514,     0.00514,
  0.00517,    0.00517,     0.00517,     0.00517,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005249,   0.005249,    0.005249,    0.005249,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004788,   0.004788,    0.004788,    0.004788,
  0.004686,   0.004686,    0.004686,    0.004686,
  0.004488,   0.004488,    0.004488,    0.004488,
  0.004309,   0.004309,    0.004309,    0.004309,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004599,   0.004599,    0.004599,    0.004599,
  0.004642,   0.004642,    0.004642,    0.004642,
  0.0047,     0.0047,      0.0047,      0.0047,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004773,   0.004773,    0.004773,    0.004773,
  0.004773,   0.004773,    0.004773,    0.004773,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004773,   0.004773,    0.004773,    0.004773,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004877,   0.004877,    0.004877,    0.004877,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004877,   0.004877,    0.004877,    0.004877,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004714,   0.004714,    0.004714,    0.004714,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004656,   0.004656,    0.004656,    0.004656,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004501,   0.004501,    0.004501,    0.004501,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004073,   0.004073,    0.004073,    0.004073,
  0.004034,   0.004034,    0.004034,    0.004034,
  0.004034,   0.004034,    0.004034,    0.004034,
  0.004047,   0.004047,    0.004047,    0.004047,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004098,   0.004098,    0.004098,    0.004098,
  0.004098,   0.004098,    0.004098,    0.004098,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004501,   0.004501,    0.004501,    0.004501,
  0.004628,   0.004628,    0.004628,    0.004628,
  0.004744,   0.004744,    0.004744,    0.004744,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004788,   0.004788,    0.004788,    0.004788,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.0047,     0.0047,      0.0047,      0.0047,
  0.004642,   0.004642,    0.004642,    0.004642,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004599,   0.004599,    0.004599,    0.004599,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004336,   0.004336,    0.004336,    0.004336,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004177,   0.004177,    0.004177,    0.004177,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.004092,   0.004092,    0.004092,    0.004092,
  0.004016,   0.004016,    0.004016,    0.004016,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.003921,   0.003921,    0.003921,    0.003921,
  0.003877,   0.003877,    0.003877,    0.003877,
  0.003883,   0.003883,    0.003883,    0.003883,
  0.003915,   0.003915,    0.003915,    0.003915,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.004034,   0.004034,    0.004034,    0.004034,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.004072,   0.004072,    0.004072,    0.004072,
  0.004072,   0.004072,    0.004072,    0.004072,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.003984,   0.003984,    0.003984,    0.003984,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.003788,   0.003788,    0.003788,    0.003788,
  0.003716,   0.003716,    0.003716,    0.003716,
  0.003716,   0.003716,    0.003716,    0.003716,
  0.003764,   0.003764,    0.003764,    0.003764,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.004098,   0.004098,    0.004098,    0.004098,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004237,   0.004237,    0.004237,    0.004237,
  0.004187,   0.004187,    0.004187,    0.004187,
  0.004156,   0.004156,    0.004156,    0.004156,
  0.004142,   0.004142,    0.004142,    0.004142,
  0.004161,   0.004161,    0.004161,    0.004161,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.004152,   0.004152,    0.004152,    0.004152,
  0.004139,   0.004139,    0.004139,    0.004139,
  0.004158,   0.004158,    0.004158,    0.004158,
  0.004137,   0.004137,    0.004137,    0.004137,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.004047,   0.004047,    0.004047,    0.004047,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.003897,   0.003897,    0.003897,    0.003897,
  0.003836,   0.003836,    0.003836,    0.003836,
  0.003788,   0.003788,    0.003788,    0.003788,
  0.003764,   0.003764,    0.003764,    0.003764,
  0.003752,   0.003752,    0.003752,    0.003752,
  0.003752,   0.003752,    0.003752,    0.003752,
  0.003776,   0.003776,    0.003776,    0.003776,
  0.003792,   0.003792,    0.003792,    0.003792,
  0.003822,   0.003822,    0.003822,    0.003822,
  0.003839,   0.003839,    0.003839,    0.003839,
  0.003845,   0.003845,    0.003845,    0.003845,
  0.003883,   0.003883,    0.003883,    0.003883,
  0.003908,   0.003908,    0.003908,    0.003908,
  0.003921,   0.003921,    0.003921,    0.003921,
  0.003954,   0.003954,    0.003954,    0.003954,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.004066,   0.004066,    0.004066,    0.004066,
  0.004102,   0.004102,    0.004102,    0.004102,
  0.004158,   0.004158,    0.004158,    0.004158,
  0.004213,   0.004213,    0.004213,    0.004213,
  0.004253,   0.004253,    0.004253,    0.004253,
  0.004293,   0.004293,    0.004293,    0.004293,
  0.004334,   0.004334,    0.004334,    0.004334,
  0.00436,    0.00436,     0.00436,     0.00436,
  0.004402,   0.004402,    0.004402,    0.004402,
  0.004478,   0.004478,    0.004478,    0.004478,
  0.00456,    0.00456,     0.00456,     0.00456,
  0.004602,   0.004602,    0.004602,    0.004602,
  0.00466,    0.00466,     0.00466,     0.00466,
  0.004755,   0.004755,    0.004755,    0.004755,
  0.004845,   0.004845,    0.004845,    0.004845,
  0.004925,   0.004925,    0.004925,    0.004925,
  0.005006,   0.005006,    0.005006,    0.005006,
  0.005089,   0.005089,    0.005089,    0.005089,
  0.005218,   0.005218,    0.005218,    0.005218,
  0.005286,   0.005286,    0.005286,    0.005286,
  0.00527,    0.00527,     0.00527,     0.00527,
  0.005333,   0.005333,    0.005333,    0.005333,
  0.005443,   0.005443,    0.005443,    0.005443,
  0.005533,   0.005533,    0.005533,    0.005533,
  0.005609,   0.005609,    0.005609,    0.005609,
  0.005672,   0.005672,    0.005672,    0.005672,
  0.005701,   0.005701,    0.005701,    0.005701,
  0.005706,   0.005706,    0.005706,    0.005706,
  0.0057,     0.0057,      0.0057,      0.0057,
  0.00569,    0.00569,     0.00569,     0.00569,
  0.005676,   0.005676,    0.005676,    0.005676,
  0.005651,   0.005651,    0.005651,    0.005651,
  0.005647,   0.005647,    0.005647,    0.005647,
  0.005718,   0.005718,    0.005718,    0.005718,
  0.005775,   0.005775,    0.005775,    0.005775,
  0.005744,   0.005744,    0.005744,    0.005744,
  0.005672,   0.005672,    0.005672,    0.005672,
  0.005561,   0.005561,    0.005561,    0.005561,
  0.005433,   0.005433,    0.005433,    0.005433,
  0.005414,   0.005414,    0.005414,    0.005414,
  0.005447,   0.005447,    0.005447,    0.005447,
  0.005349,   0.005349,    0.005349,    0.005349,
  0.005186,   0.005186,    0.005186,    0.005186,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005202,   0.005202,    0.005202,    0.005202,
  0.005202,   0.005202,    0.005202,    0.005202,
  0.005219,   0.005219,    0.005219,    0.005219,
  0.005269,   0.005269,    0.005269,    0.005269,
  0.005334,   0.005334,    0.005334,    0.005334,
  0.005353,   0.005353,    0.005353,    0.005353,
  0.005405,   0.005405,    0.005405,    0.005405,
  0.00548,    0.00548,     0.00548,     0.00548,
  0.005525,   0.005525,    0.005525,    0.005525,
  0.005564,   0.005564,    0.005564,    0.005564,
  0.005586,   0.005586,    0.005586,    0.005586,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005564,   0.005564,    0.005564,    0.005564,
  0.005511,   0.005511,    0.005511,    0.005511,
  0.00547,    0.00547,     0.00547,     0.00547,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.005327,   0.005327,    0.005327,    0.005327,
  0.005237,   0.005237,    0.005237,    0.005237,
  0.005171,   0.005171,    0.005171,    0.005171,
  0.005045,   0.005045,    0.005045,    0.005045,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004628,   0.004628,    0.004628,    0.004628,
  0.004744,   0.004744,    0.004744,    0.004744,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004803,   0.004803,    0.004803,    0.004803,
  0.004953,   0.004953,    0.004953,    0.004953,
  0.004953,   0.004953,    0.004953,    0.004953,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004967,   0.004967,    0.004967,    0.004967,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004788,   0.004788,    0.004788,    0.004788,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004686,   0.004686,    0.004686,    0.004686,
  0.004657,   0.004657,    0.004657,    0.004657,
  0.004818,   0.004818,    0.004818,    0.004818,
  0.005045,   0.005045,    0.005045,    0.005045,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005266,   0.005266,    0.005266,    0.005266,
  0.005478,   0.005478,    0.005478,    0.005478,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005562,   0.005562,    0.005562,    0.005562,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005494,   0.005494,    0.005494,    0.005494,
  0.005174,   0.005174,    0.005174,    0.005174,
  0.004833,   0.004833,    0.004833,    0.004833,
  0.004519,   0.004519,    0.004519,    0.004519,
  0.004216,   0.004216,    0.004216,    0.004216,
  0.004023,   0.004023,    0.004023,    0.004023,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003872,   0.003872,    0.003872,    0.003872,
  0.003776,   0.003776,    0.003776,    0.003776,
  0.003669,   0.003669,    0.003669,    0.003669,
  0.003646,   0.003646,    0.003646,    0.003646,
  0.003646,   0.003646,    0.003646,    0.003646,
  0.003623,   0.003623,    0.003623,    0.003623,
  0.003577,   0.003577,    0.003577,    0.003577,
  0.00352,    0.00352,     0.00352,     0.00352,
  0.003509,   0.003509,    0.003509,    0.003509,
  0.003465,   0.003465,    0.003465,    0.003465,
  0.003377,   0.003377,    0.003377,    0.003377,
  0.003377,   0.003377,    0.003377,    0.003377,
  0.003377,   0.003377,    0.003377,    0.003377,
  0.003355,   0.003355,    0.003355,    0.003355,
  0.003334,   0.003334,    0.003334,    0.003334,
  0.003323,   0.003323,    0.003323,    0.003323,
  0.003334,   0.003334,    0.003334,    0.003334,
  0.003291,   0.003291,    0.003291,    0.003291,
  0.00327,    0.00327,     0.00327,     0.00327,
  0.003281,   0.003281,    0.003281,    0.003281,
  0.003323,   0.003323,    0.003323,    0.003323,
  0.003302,   0.003302,    0.003302,    0.003302,
  0.003228,   0.003228,    0.003228,    0.003228,
  0.003239,   0.003239,    0.003239,    0.003239,
  0.003239,   0.003239,    0.003239,    0.003239,
  0.003239,   0.003239,    0.003239,    0.003239,
  0.003281,   0.003281,    0.003281,    0.003281,
  0.003367,   0.003367,    0.003367,    0.003367,
  0.003465,   0.003465,    0.003465,    0.003465,
  0.003601,   0.003601,    0.003601,    0.003601,
  0.003838,   0.003838,    0.003838,    0.003838,
  0.004181,   0.004181,    0.004181,    0.004181,
  0.004603,   0.004603,    0.004603,    0.004603,
  0.004954,   0.004954,    0.004954,    0.004954,
  0.005016,   0.005016,    0.005016,    0.005016,
  0.004889,   0.004889,    0.004889,    0.004889,
  0.004926,   0.004926,    0.004926,    0.004926,
  0.004997,   0.004997,    0.004997,    0.004997,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.00477,    0.00477,     0.00477,     0.00477,
  0.004483,   0.004483,    0.004483,    0.004483,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004212,   0.004212,    0.004212,    0.004212,
  0.004098,   0.004098,    0.004098,    0.004098,
  0.003869,   0.003869,    0.003869,    0.003869,
  0.00367,    0.00367,     0.00367,     0.00367,
  0.003577,   0.003577,    0.003577,    0.003577,
  0.003577,   0.003577,    0.003577,    0.003577,
  0.003566,   0.003566,    0.003566,    0.003566,
  0.003566,   0.003566,    0.003566,    0.003566,
  0.003611,   0.003611,    0.003611,    0.003611,
  0.003646,   0.003646,    0.003646,    0.003646,
  0.003658,   0.003658,    0.003658,    0.003658,
  0.003658,   0.003658,    0.003658,    0.003658,
  0.003669,   0.003669,    0.003669,    0.003669,
  0.003693,   0.003693,    0.003693,    0.003693,
  0.003704,   0.003704,    0.003704,    0.003704,
  0.003693,   0.003693,    0.003693,    0.003693,
  0.003693,   0.003693,    0.003693,    0.003693,
  0.00374,    0.00374,     0.00374,     0.00374,
  0.003788,   0.003788,    0.003788,    0.003788,
  0.0038,     0.0038,      0.0038,      0.0038,
  0.0038,     0.0038,      0.0038,      0.0038,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.0038,     0.0038,      0.0038,      0.0038,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.003836,   0.003836,    0.003836,    0.003836,
  0.00386,    0.00386,     0.00386,     0.00386,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.003922,   0.003922,    0.003922,    0.003922,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003897,   0.003897,    0.003897,    0.003897,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.003872,   0.003872,    0.003872,    0.003872,
  0.003872,   0.003872,    0.003872,    0.003872,
  0.00386,    0.00386,     0.00386,     0.00386,
  0.003848,   0.003848,    0.003848,    0.003848,
  0.003848,   0.003848,    0.003848,    0.003848,
  0.00386,    0.00386,     0.00386,     0.00386,
  0.003848,   0.003848,    0.003848,    0.003848,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.003776,   0.003776,    0.003776,    0.003776,
  0.003728,   0.003728,    0.003728,    0.003728,
  0.003681,   0.003681,    0.003681,    0.003681,
  0.003646,   0.003646,    0.003646,    0.003646,
  0.003634,   0.003634,    0.003634,    0.003634,
  0.003623,   0.003623,    0.003623,    0.003623,
  0.003623,   0.003623,    0.003623,    0.003623,
  0.0036,     0.0036,      0.0036,      0.0036,
  0.003532,   0.003532,    0.003532,    0.003532,
  0.003465,   0.003465,    0.003465,    0.003465,
  0.00341,    0.00341,     0.00341,     0.00341,
  0.003355,   0.003355,    0.003355,    0.003355,
  0.003302,   0.003302,    0.003302,    0.003302,
  0.003281,   0.003281,    0.003281,    0.003281,
  0.003249,   0.003249,    0.003249,    0.003249,
  0.003197,   0.003197,    0.003197,    0.003197,
  0.003146,   0.003146,    0.003146,    0.003146,
  0.003095,   0.003095,    0.003095,    0.003095,
  0.003055,   0.003055,    0.003055,    0.003055,
  0.003016,   0.003016,    0.003016,    0.003016,
  0.002987,   0.002987,    0.002987,    0.002987,
  0.002967,   0.002967,    0.002967,    0.002967,
  0.002948,   0.002948,    0.002948,    0.002948,
  0.002919,   0.002919,    0.002919,    0.002919,
  0.002881,   0.002881,    0.002881,    0.002881,
  0.002881,   0.002881,    0.002881,    0.002881,
  0.002919,   0.002919,    0.002919,    0.002919,
  0.002938,   0.002938,    0.002938,    0.002938,
  0.002929,   0.002929,    0.002929,    0.002929,
  0.002919,   0.002919,    0.002919,    0.002919,
  0.00291,    0.00291,     0.00291,     0.00291,
  0.002881,   0.002881,    0.002881,    0.002881,
  0.002835,   0.002835,    0.002835,    0.002835,
  0.002798,   0.002798,    0.002798,    0.002798,
  0.00277,    0.00277,     0.00277,     0.00277,
  0.002716,   0.002716,    0.002716,    0.002716,
  0.002707,   0.002707,    0.002707,    0.002707,
  0.002761,   0.002761,    0.002761,    0.002761,
  0.002798,   0.002798,    0.002798,    0.002798,
  0.002863,   0.002863,    0.002863,    0.002863,
  0.002977,   0.002977,    0.002977,    0.002977,
  0.003096,   0.003096,    0.003096,    0.003096,
  0.003197,   0.003197,    0.003197,    0.003197,
  0.003281,   0.003281,    0.003281,    0.003281,
  0.003377,   0.003377,    0.003377,    0.003377,
  0.003431,   0.003431,    0.003431,    0.003431,
  0.003454,   0.003454,    0.003454,    0.003454,
  0.003498,   0.003498,    0.003498,    0.003498,
  0.00352,    0.00352,     0.00352,     0.00352,
  0.00352,    0.00352,     0.00352,     0.00352,
  0.00352,    0.00352,     0.00352,     0.00352,
  0.00352,    0.00352,     0.00352,     0.00352,
  0.003498,   0.003498,    0.003498,    0.003498,
  0.003443,   0.003443,    0.003443,    0.003443,
  0.00341,    0.00341,     0.00341,     0.00341,
  0.003399,   0.003399,    0.003399,    0.003399,
  0.003377,   0.003377,    0.003377,    0.003377,
  0.003334,   0.003334,    0.003334,    0.003334,
  0.003312,   0.003312,    0.003312,    0.003312,
  0.003291,   0.003291,    0.003291,    0.003291,
  0.003218,   0.003218,    0.003218,    0.003218,
  0.003116,   0.003116,    0.003116,    0.003116,
  0.003075,   0.003075,    0.003075,    0.003075,
  0.003146,   0.003146,    0.003146,    0.003146,
  0.003156,   0.003156,    0.003156,    0.003156,
  0.003056,   0.003056,    0.003056,    0.003056,
  0.002977,   0.002977,    0.002977,    0.002977,
  0.002987,   0.002987,    0.002987,    0.002987,
  0.003036,   0.003036,    0.003036,    0.003036,
  0.003085,   0.003085,    0.003085,    0.003085,
  0.003146,   0.003146,    0.003146,    0.003146,
  0.003207,   0.003207,    0.003207,    0.003207,
  0.00327,    0.00327,     0.00327,     0.00327,
  0.003345,   0.003345,    0.003345,    0.003345,
  0.00341,    0.00341,     0.00341,     0.00341,
  0.003454,   0.003454,    0.003454,    0.003454,
  0.003476,   0.003476,    0.003476,    0.003476,
  0.003532,   0.003532,    0.003532,    0.003532,
  0.003611,   0.003611,    0.003611,    0.003611,
  0.003669,   0.003669,    0.003669,    0.003669,
  0.003728,   0.003728,    0.003728,    0.003728,
  0.003788,   0.003788,    0.003788,    0.003788,
  0.003848,   0.003848,    0.003848,    0.003848,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.003897,   0.003897,    0.003897,    0.003897,
  0.003922,   0.003922,    0.003922,    0.003922,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.004176,   0.004176,    0.004176,    0.004176,
  0.004296,   0.004296,    0.004296,    0.004296,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004585,   0.004585,    0.004585,    0.004585,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004585,   0.004585,    0.004585,    0.004585,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004336,   0.004336,    0.004336,    0.004336,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004176,   0.004176,    0.004176,    0.004176,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004309,   0.004309,    0.004309,    0.004309,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004137,   0.004137,    0.004137,    0.004137,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004072,   0.004072,    0.004072,    0.004072,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004472,   0.004472,    0.004472,    0.004472,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004585,   0.004585,    0.004585,    0.004585,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004308,   0.004308,    0.004308,    0.004308,
  0.004308,   0.004308,    0.004308,    0.004308,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.003897,   0.003897,    0.003897,    0.003897,
  0.003836,   0.003836,    0.003836,    0.003836,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.0047,     0.0047,      0.0047,      0.0047,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004771,   0.004771,    0.004771,    0.004771,
  0.004635,   0.004635,    0.004635,    0.004635,
  0.004453,   0.004453,    0.004453,    0.004453,
  0.004333,   0.004333,    0.004333,    0.004333,
  0.004276,   0.004276,    0.004276,    0.004276,
  0.00427,    0.00427,     0.00427,     0.00427,
  0.004278,   0.004278,    0.004278,    0.004278,
  0.004232,   0.004232,    0.004232,    0.004232,
  0.004138,   0.004138,    0.004138,    0.004138,
  0.004061,   0.004061,    0.004061,    0.004061,
  0.004016,   0.004016,    0.004016,    0.004016,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.003908,   0.003908,    0.003908,    0.003908,
  0.003845,   0.003845,    0.003845,    0.003845,
  0.003818,   0.003818,    0.003818,    0.003818,
  0.003791,   0.003791,    0.003791,    0.003791,
  0.003746,   0.003746,    0.003746,    0.003746,
  0.003751,   0.003751,    0.003751,    0.003751,
  0.003787,   0.003787,    0.003787,    0.003787,
  0.003798,   0.003798,    0.003798,    0.003798,
  0.00374,    0.00374,     0.00374,     0.00374,
  0.00363,    0.00363,     0.00363,     0.00363,
  0.003599,   0.003599,    0.003599,    0.003599,
  0.003591,   0.003591,    0.003591,    0.003591,
  0.003541,   0.003541,    0.003541,    0.003541,
  0.003491,   0.003491,    0.003491,    0.003491,
  0.003423,   0.003423,    0.003423,    0.003423,
  0.00336,    0.00336,     0.00336,     0.00336,
  0.003383,   0.003383,    0.003383,    0.003383,
  0.00337,    0.00337,     0.00337,     0.00337,
  0.003357,   0.003357,    0.003357,    0.003357,
  0.003362,   0.003362,    0.003362,    0.003362,
  0.003318,   0.003318,    0.003318,    0.003318,
  0.003318,   0.003318,    0.003318,    0.003318,
  0.003318,   0.003318,    0.003318,    0.003318,
  0.003318,   0.003318,    0.003318,    0.003318,
  0.00337,    0.00337,     0.00337,     0.00337,
  0.00336,    0.00336,     0.00336,     0.00336,
  0.003211,   0.003211,    0.003211,    0.003211,
  0.003093,   0.003093,    0.003093,    0.003093,
  0.003103,   0.003103,    0.003103,    0.003103,
  0.00313,    0.00313,     0.00313,     0.00313,
  0.003112,   0.003112,    0.003112,    0.003112,
  0.003063,   0.003063,    0.003063,    0.003063,
  0.003045,   0.003045,    0.003045,    0.003045,
  0.003031,   0.003031,    0.003031,    0.003031,
  0.003035,   0.003035,    0.003035,    0.003035,
  0.003071,   0.003071,    0.003071,    0.003071,
  0.003093,   0.003093,    0.003093,    0.003093,
  0.003116,   0.003116,    0.003116,    0.003116,
  0.003139,   0.003139,    0.003139,    0.003139,
  0.003131,   0.003131,    0.003131,    0.003131,
  0.003129,   0.003129,    0.003129,    0.003129,
  0.003153,   0.003153,    0.003153,    0.003153,
  0.003203,   0.003203,    0.003203,    0.003203,
  0.003234,   0.003234,    0.003234,    0.003234,
  0.003215,   0.003215,    0.003215,    0.003215,
  0.003204,   0.003204,    0.003204,    0.003204,
  0.003185,   0.003185,    0.003185,    0.003185,
  0.003194,   0.003194,    0.003194,    0.003194,
  0.003208,   0.003208,    0.003208,    0.003208,
  0.003217,   0.003217,    0.003217,    0.003217,
  0.003196,   0.003196,    0.003196,    0.003196,
  0.003154,   0.003154,    0.003154,    0.003154,
  0.003163,   0.003163,    0.003163,    0.003163,
  0.003161,   0.003161,    0.003161,    0.003161,
  0.003138,   0.003138,    0.003138,    0.003138,
  0.003148,   0.003148,    0.003148,    0.003148,
  0.003158,   0.003158,    0.003158,    0.003158,
  0.003158,   0.003158,    0.003158,    0.003158,
  0.003156,   0.003156,    0.003156,    0.003156,
  0.003166,   0.003166,    0.003166,    0.003166,
  0.003165,   0.003165,    0.003165,    0.003165,
  0.003144,   0.003144,    0.003144,    0.003144,
  0.003123,   0.003123,    0.003123,    0.003123,
  0.003134,   0.003134,    0.003134,    0.003134,
  0.003144,   0.003144,    0.003144,    0.003144,
  0.003155,   0.003155,    0.003155,    0.003155,
  0.003165,   0.003165,    0.003165,    0.003165,
  0.003165,   0.003165,    0.003165,    0.003165,
  0.003176,   0.003176,    0.003176,    0.003176,
  0.003186,   0.003186,    0.003186,    0.003186,
  0.003229,   0.003229,    0.003229,    0.003229,
  0.003299,   0.003299,    0.003299,    0.003299,
  0.003335,   0.003335,    0.003335,    0.003335,
  0.003395,   0.003395,    0.003395,    0.003395,
  0.003436,   0.003436,    0.003436,    0.003436,
  0.00343,    0.00343,     0.00343,     0.00343,
  0.003437,   0.003437,    0.003437,    0.003437,
  0.003478,   0.003478,    0.003478,    0.003478,
  0.003557,   0.003557,    0.003557,    0.003557,
  0.003597,   0.003597,    0.003597,    0.003597,
  0.003656,   0.003656,    0.003656,    0.003656,
  0.003669,   0.003669,    0.003669,    0.003669,
  0.003645,   0.003645,    0.003645,    0.003645,
  0.003678,   0.003678,    0.003678,    0.003678,
  0.003698,   0.003698,    0.003698,    0.003698,
  0.003717,   0.003717,    0.003717,    0.003717,
  0.003749,   0.003749,    0.003749,    0.003749,
  0.00378,    0.00378,     0.00378,     0.00378,
  0.0038,     0.0038,      0.0038,      0.0038,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.003824,   0.003824,    0.003824,    0.003824,
  0.003836,   0.003836,    0.003836,    0.003836,
  0.00386,    0.00386,     0.00386,     0.00386,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.003897,   0.003897,    0.003897,    0.003897,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003922,   0.003922,    0.003922,    0.003922,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.003984,   0.003984,    0.003984,    0.003984,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.004034,   0.004034,    0.004034,    0.004034,
  0.003984,   0.003984,    0.003984,    0.003984,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003897,   0.003897,    0.003897,    0.003897,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004098,   0.004098,    0.004098,    0.004098,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004137,   0.004137,    0.004137,    0.004137,
  0.004047,   0.004047,    0.004047,    0.004047,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.004034,   0.004034,    0.004034,    0.004034,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004137,   0.004137,    0.004137,    0.004137,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004137,   0.004137,    0.004137,    0.004137,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004047,   0.004047,    0.004047,    0.004047,
  0.004047,   0.004047,    0.004047,    0.004047,
  0.004047,   0.004047,    0.004047,    0.004047,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.004047,   0.004047,    0.004047,    0.004047,
  0.004098,   0.004098,    0.004098,    0.004098,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.004073,   0.004073,    0.004073,    0.004073,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003922,   0.003922,    0.003922,    0.003922,
  0.00389,    0.00389,     0.00389,     0.00389,
  0.003859,   0.003859,    0.003859,    0.003859,
  0.003839,   0.003839,    0.003839,    0.003839,
  0.003845,   0.003845,    0.003845,    0.003845,
  0.003896,   0.003896,    0.003896,    0.003896,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.004037,   0.004037,    0.004037,    0.004037,
  0.004084,   0.004084,    0.004084,    0.004084,
  0.00412,    0.00412,     0.00412,     0.00412,
  0.004174,   0.004174,    0.004174,    0.004174,
  0.004201,   0.004201,    0.004201,    0.004201,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004266,   0.004266,    0.004266,    0.004266,
  0.004302,   0.004302,    0.004302,    0.004302,
  0.004356,   0.004356,    0.004356,    0.004356,
  0.004414,   0.004414,    0.004414,    0.004414,
  0.004471,   0.004471,    0.004471,    0.004471,
  0.004513,   0.004513,    0.004513,    0.004513,
  0.00451,    0.00451,     0.00451,     0.00451,
  0.004541,   0.004541,    0.004541,    0.004541,
  0.004603,   0.004603,    0.004603,    0.004603,
  0.00465,    0.00465,     0.00465,     0.00465,
  0.004744,   0.004744,    0.004744,    0.004744,
  0.00487,    0.00487,     0.00487,     0.00487,
  0.004965,   0.004965,    0.004965,    0.004965,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005218,   0.005218,    0.005218,    0.005218,
  0.005298,   0.005298,    0.005298,    0.005298,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005444,   0.005444,    0.005444,    0.005444,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005269,   0.005269,    0.005269,    0.005269,
  0.004864,   0.004864,    0.004864,    0.004864,
  0.004671,   0.004671,    0.004671,    0.004671,
  0.004642,   0.004642,    0.004642,    0.004642,
  0.004628,   0.004628,    0.004628,    0.004628,
  0.004599,   0.004599,    0.004599,    0.004599,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004544,   0.004544,    0.004544,    0.004544,
  0.004711,   0.004711,    0.004711,    0.004711,
  0.004795,   0.004795,    0.004795,    0.004795,
  0.004855,   0.004855,    0.004855,    0.004855,
  0.004871,   0.004871,    0.004871,    0.004871,
  0.004794,   0.004794,    0.004794,    0.004794,
  0.004639,   0.004639,    0.004639,    0.004639,
  0.004623,   0.004623,    0.004623,    0.004623,
  0.004715,   0.004715,    0.004715,    0.004715,
  0.004777,   0.004777,    0.004777,    0.004777,
  0.004794,   0.004794,    0.004794,    0.004794,
  0.004793,   0.004793,    0.004793,    0.004793,
  0.004855,   0.004855,    0.004855,    0.004855,
  0.004902,   0.004902,    0.004902,    0.004902,
  0.004871,   0.004871,    0.004871,    0.004871,
  0.004734,   0.004734,    0.004734,    0.004734,
  0.004541,   0.004541,    0.004541,    0.004541,
  0.004382,   0.004382,    0.004382,    0.004382,
  0.00427,    0.00427,     0.00427,     0.00427,
  0.00426,    0.00426,     0.00426,     0.00426,
  0.004305,   0.004305,    0.004305,    0.004305,
  0.004296,   0.004296,    0.004296,    0.004296,
  0.004237,   0.004237,    0.004237,    0.004237,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.004098,   0.004098,    0.004098,    0.004098,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004072,   0.004072,    0.004072,    0.004072,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004176,   0.004176,    0.004176,    0.004176,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004308,   0.004308,    0.004308,    0.004308,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004473,   0.004473,    0.004473,    0.004473,
  0.0046,     0.0046,      0.0046,      0.0046,
  0.004789,   0.004789,    0.004789,    0.004789,
  0.004951,   0.004951,    0.004951,    0.004951,
  0.004999,   0.004999,    0.004999,    0.004999,
  0.004995,   0.004995,    0.004995,    0.004995,
  0.004979,   0.004979,    0.004979,    0.004979,
  0.004962,   0.004962,    0.004962,    0.004962,
  0.00497,    0.00497,     0.00497,     0.00497,
  0.004956,   0.004956,    0.004956,    0.004956,
  0.004961,   0.004961,    0.004961,    0.004961,
  0.005015,   0.005015,    0.005015,    0.005015,
  0.005002,   0.005002,    0.005002,    0.005002,
  0.004939,   0.004939,    0.004939,    0.004939,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004808,   0.004808,    0.004808,    0.004808,
  0.004641,   0.004641,    0.004641,    0.004641,
  0.004584,   0.004584,    0.004584,    0.004584,
  0.004555,   0.004555,    0.004555,    0.004555,
  0.004446,   0.004446,    0.004446,    0.004446,
  0.004232,   0.004232,    0.004232,    0.004232,
  0.004039,   0.004039,    0.004039,    0.004039,
  0.003926,   0.003926,    0.003926,    0.003926,
  0.003831,   0.003831,    0.003831,    0.003831,
  0.003768,   0.003768,    0.003768,    0.003768,
  0.003704,   0.003704,    0.003704,    0.003704,
  0.003673,   0.003673,    0.003673,    0.003673,
  0.003704,   0.003704,    0.003704,    0.003704,
  0.003815,   0.003815,    0.003815,    0.003815,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003957,   0.003957,    0.003957,    0.003957,
  0.00402,    0.00402,     0.00402,     0.00402,
  0.004068,   0.004068,    0.004068,    0.004068,
  0.004083,   0.004083,    0.004083,    0.004083,
  0.004083,   0.004083,    0.004083,    0.004083,
  0.004067,   0.004067,    0.004067,    0.004067,
  0.004051,   0.004051,    0.004051,    0.004051,
  0.004067,   0.004067,    0.004067,    0.004067,
  0.004067,   0.004067,    0.004067,    0.004067,
  0.004052,   0.004052,    0.004052,    0.004052,
  0.004052,   0.004052,    0.004052,    0.004052,
  0.004068,   0.004068,    0.004068,    0.004068,
  0.0041,     0.0041,      0.0041,      0.0041,
  0.004147,   0.004147,    0.004147,    0.004147,
  0.004336,   0.004336,    0.004336,    0.004336,
  0.004636,   0.004636,    0.004636,    0.004636,
  0.004781,   0.004781,    0.004781,    0.004781,
  0.004682,   0.004682,    0.004682,    0.004682,
  0.004555,   0.004555,    0.004555,    0.004555,
  0.004601,   0.004601,    0.004601,    0.004601,
  0.004659,   0.004659,    0.004659,    0.004659,
  0.004737,   0.004737,    0.004737,    0.004737,
  0.004965,   0.004965,    0.004965,    0.004965,
  0.005171,   0.005171,    0.005171,    0.005171,
  0.005234,   0.005234,    0.005234,    0.005234,
  0.005218,   0.005218,    0.005218,    0.005218,
  0.005191,   0.005191,    0.005191,    0.005191,
  0.005183,   0.005183,    0.005183,    0.005183,
  0.005227,   0.005227,    0.005227,    0.005227,
  0.005278,   0.005278,    0.005278,    0.005278,
  0.005317,   0.005317,    0.005317,    0.005317,
  0.005348,   0.005348,    0.005348,    0.005348,
  0.005554,   0.005554,    0.005554,    0.005554,
  0.005823,   0.005823,    0.005823,    0.005823,
  0.00591,    0.00591,     0.00591,     0.00591,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.005766,   0.005766,    0.005766,    0.005766,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005186,   0.005186,    0.005186,    0.005186,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.004848,   0.004848,    0.004848,    0.004848,
  0.004671,   0.004671,    0.004671,    0.004671,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004112,   0.004112,    0.004112,    0.004112,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.00386,    0.00386,     0.00386,     0.00386,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.003788,   0.003788,    0.003788,    0.003788,
  0.003788,   0.003788,    0.003788,    0.003788,
  0.003752,   0.003752,    0.003752,    0.003752,
  0.003669,   0.003669,    0.003669,    0.003669,
  0.003646,   0.003646,    0.003646,    0.003646,
  0.003634,   0.003634,    0.003634,    0.003634,
  0.0036,     0.0036,      0.0036,      0.0036,
  0.0036,     0.0036,      0.0036,      0.0036,
  0.003634,   0.003634,    0.003634,    0.003634,
  0.003693,   0.003693,    0.003693,    0.003693,
  0.003752,   0.003752,    0.003752,    0.003752,
  0.003776,   0.003776,    0.003776,    0.003776,
  0.003836,   0.003836,    0.003836,    0.003836,
  0.004049,   0.004049,    0.004049,    0.004049,
  0.00431,    0.00431,     0.00431,     0.00431,
  0.004632,   0.004632,    0.004632,    0.004632,
  0.005,      0.005,       0.005,       0.005,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005132,   0.005132,    0.005132,    0.005132,
  0.004924,   0.004924,    0.004924,    0.004924,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004869,   0.004869,    0.004869,    0.004869,
  0.004889,   0.004889,    0.004889,    0.004889,
  0.004886,   0.004886,    0.004886,    0.004886,
  0.004872,   0.004872,    0.004872,    0.004872,
  0.004814,   0.004814,    0.004814,    0.004814,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.0046,     0.0046,      0.0046,      0.0046,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004501,   0.004501,    0.004501,    0.004501,
  0.004686,   0.004686,    0.004686,    0.004686,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.00551,    0.00551,     0.00551,     0.00551,
  0.005445,   0.005445,    0.005445,    0.005445,
  0.005366,   0.005366,    0.005366,    0.005366,
  0.005301,   0.005301,    0.005301,    0.005301,
  0.005238,   0.005238,    0.005238,    0.005238,
  0.00519,    0.00519,     0.00519,     0.00519,
  0.005172,   0.005172,    0.005172,    0.005172,
  0.005123,   0.005123,    0.005123,    0.005123,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.00538,    0.00538,     0.00538,     0.00538,
  0.005524,   0.005524,    0.005524,    0.005524,
  0.005664,   0.005664,    0.005664,    0.005664,
  0.005788,   0.005788,    0.005788,    0.005788,
  0.005968,   0.005968,    0.005968,    0.005968,
  0.00612,    0.00612,     0.00612,     0.00612,
  0.006153,   0.006153,    0.006153,    0.006153,
  0.006171,   0.006171,    0.006171,    0.006171,
  0.00611,    0.00611,     0.00611,     0.00611,
  0.005947,   0.005947,    0.005947,    0.005947,
  0.005842,   0.005842,    0.005842,    0.005842,
  0.005822,   0.005822,    0.005822,    0.005822,
  0.005856,   0.005856,    0.005856,    0.005856,
  0.005984,   0.005984,    0.005984,    0.005984,
  0.006131,   0.006131,    0.006131,    0.006131,
  0.006151,   0.006151,    0.006151,    0.006151,
  0.006162,   0.006162,    0.006162,    0.006162,
  0.006176,   0.006176,    0.006176,    0.006176,
  0.006179,   0.006179,    0.006179,    0.006179,
  0.006171,   0.006171,    0.006171,    0.006171,
  0.006136,   0.006136,    0.006136,    0.006136,
  0.00609,    0.00609,     0.00609,     0.00609,
  0.005988,   0.005988,    0.005988,    0.005988,
  0.005894,   0.005894,    0.005894,    0.005894,
  0.005799,   0.005799,    0.005799,    0.005799,
  0.005729,   0.005729,    0.005729,    0.005729,
  0.005635,   0.005635,    0.005635,    0.005635,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.005497,   0.005497,    0.005497,    0.005497,
  0.00561,    0.00561,     0.00561,     0.00561,
  0.005773,   0.005773,    0.005773,    0.005773,
  0.005868,   0.005868,    0.005868,    0.005868,
  0.005837,   0.005837,    0.005837,    0.005837,
  0.005732,   0.005732,    0.005732,    0.005732,
  0.005614,   0.005614,    0.005614,    0.005614,
  0.005551,   0.005551,    0.005551,    0.005551,
  0.005533,   0.005533,    0.005533,    0.005533,
  0.00551,    0.00551,     0.00551,     0.00551,
  0.005452,   0.005452,    0.005452,    0.005452,
  0.005409,   0.005409,    0.005409,    0.005409,
  0.005388,   0.005388,    0.005388,    0.005388,
  0.005302,   0.005302,    0.005302,    0.005302,
  0.005199,   0.005199,    0.005199,    0.005199,
  0.005151,   0.005151,    0.005151,    0.005151,
  0.005139,   0.005139,    0.005139,    0.005139,
  0.005158,   0.005158,    0.005158,    0.005158,
  0.005178,   0.005178,    0.005178,    0.005178,
  0.005188,   0.005188,    0.005188,    0.005188,
  0.005218,   0.005218,    0.005218,    0.005218,
  0.005213,   0.005213,    0.005213,    0.005213,
  0.005241,   0.005241,    0.005241,    0.005241,
  0.005315,   0.005315,    0.005315,    0.005315,
  0.005358,   0.005358,    0.005358,    0.005358,
  0.005401,   0.005401,    0.005401,    0.005401,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.005421,   0.005421,    0.005421,    0.005421,
  0.005377,   0.005377,    0.005377,    0.005377,
  0.005346,   0.005346,    0.005346,    0.005346,
  0.005453,   0.005453,    0.005453,    0.005453,
  0.005629,   0.005629,    0.005629,    0.005629,
  0.005862,   0.005862,    0.005862,    0.005862,
  0.006107,   0.006107,    0.006107,    0.006107,
  0.00624,    0.00624,     0.00624,     0.00624,
  0.006322,   0.006322,    0.006322,    0.006322,
  0.006436,   0.006436,    0.006436,    0.006436,
  0.006557,   0.006557,    0.006557,    0.006557,
  0.006584,   0.006584,    0.006584,    0.006584,
  0.006129,   0.006129,    0.006129,    0.006129,
  0.005499,   0.005499,    0.005499,    0.005499,
  0.005177,   0.005177,    0.005177,    0.005177,
  0.004954,   0.004954,    0.004954,    0.004954,
  0.004752,   0.004752,    0.004752,    0.004752,
  0.00454,    0.00454,     0.00454,     0.00454,
  0.00433,    0.00433,     0.00433,     0.00433,
  0.004199,   0.004199,    0.004199,    0.004199,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.00369,    0.00369,     0.00369,     0.00369,
  0.003517,   0.003517,    0.003517,    0.003517,
  0.003532,   0.003532,    0.003532,    0.003532,
  0.003563,   0.003563,    0.003563,    0.003563,
  0.00361,    0.00361,     0.00361,     0.00361,
  0.003626,   0.003626,    0.003626,    0.003626,
  0.003626,   0.003626,    0.003626,    0.003626,
  0.003693,   0.003693,    0.003693,    0.003693,
  0.003795,   0.003795,    0.003795,    0.003795,
  0.003852,   0.003852,    0.003852,    0.003852,
  0.003857,   0.003857,    0.003857,    0.003857,
  0.003855,   0.003855,    0.003855,    0.003855,
  0.003866,   0.003866,    0.003866,    0.003866,
  0.003898,   0.003898,    0.003898,    0.003898,
  0.003935,   0.003935,    0.003935,    0.003935,
  0.004018,   0.004018,    0.004018,    0.004018,
  0.004141,   0.004141,    0.004141,    0.004141,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004264,   0.004264,    0.004264,    0.004264,
  0.00432,    0.00432,     0.00432,     0.00432,
  0.004414,   0.004414,    0.004414,    0.004414,
  0.004497,   0.004497,    0.004497,    0.004497,
  0.004556,   0.004556,    0.004556,    0.004556,
  0.004622,   0.004622,    0.004622,    0.004622,
  0.004741,   0.004741,    0.004741,    0.004741,
  0.004849,   0.004849,    0.004849,    0.004849,
  0.004826,   0.004826,    0.004826,    0.004826,
  0.004769,   0.004769,    0.004769,    0.004769,
  0.004735,   0.004735,    0.004735,    0.004735,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004661,   0.004661,    0.004661,    0.004661,
  0.004624,   0.004624,    0.004624,    0.004624,
  0.004574,   0.004574,    0.004574,    0.004574,
  0.004525,   0.004525,    0.004525,    0.004525,
  0.004506,   0.004506,    0.004506,    0.004506,
  0.004497,   0.004497,    0.004497,    0.004497,
  0.00444,    0.00444,     0.00444,     0.00444,
  0.004401,   0.004401,    0.004401,    0.004401,
  0.004408,   0.004408,    0.004408,    0.004408,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004477,   0.004477,    0.004477,    0.004477,
  0.004606,   0.004606,    0.004606,    0.004606,
  0.004689,   0.004689,    0.004689,    0.004689,
  0.004706,   0.004706,    0.004706,    0.004706,
  0.004732,   0.004732,    0.004732,    0.004732,
  0.004851,   0.004851,    0.004851,    0.004851,
  0.005018,   0.005018,    0.005018,    0.005018,
  0.005108,   0.005108,    0.005108,    0.005108,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005249,   0.005249,    0.005249,    0.005249,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005646,   0.005646,    0.005646,    0.005646,
  0.005854,   0.005854,    0.005854,    0.005854,
  0.006106,   0.006106,    0.006106,    0.006106,
  0.006424,   0.006424,    0.006424,    0.006424,
  0.006716,   0.006716,    0.006716,    0.006716,
  0.006876,   0.006876,    0.006876,    0.006876,
  0.006864,   0.006864,    0.006864,    0.006864,
  0.006833,   0.006833,    0.006833,    0.006833,
  0.006804,   0.006804,    0.006804,    0.006804,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006683,   0.006683,    0.006683,    0.006683,
  0.006644,   0.006644,    0.006644,    0.006644,
  0.006616,   0.006616,    0.006616,    0.006616,
  0.006577,   0.006577,    0.006577,    0.006577,
  0.006577,   0.006577,    0.006577,    0.006577,
  0.006636,   0.006636,    0.006636,    0.006636,
  0.006675,   0.006675,    0.006675,    0.006675,
  0.006655,   0.006655,    0.006655,    0.006655,
  0.006636,   0.006636,    0.006636,    0.006636,
  0.006675,   0.006675,    0.006675,    0.006675,
  0.006775,   0.006775,    0.006775,    0.006775,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006916,   0.006916,    0.006916,    0.006916,
  0.006978,   0.006978,    0.006978,    0.006978,
  0.006987,   0.006987,    0.006987,    0.006987,
  0.006966,   0.006966,    0.006966,    0.006966,
  0.006937,   0.006937,    0.006937,    0.006937,
  0.006937,   0.006937,    0.006937,    0.006937,
  0.006966,   0.006966,    0.006966,    0.006966,
  0.006934,   0.006934,    0.006934,    0.006934,
  0.006934,   0.006934,    0.006934,    0.006934,
  0.006924,   0.006924,    0.006924,    0.006924,
  0.006935,   0.006935,    0.006935,    0.006935,
  0.006937,   0.006937,    0.006937,    0.006937,
  0.006875,   0.006875,    0.006875,    0.006875,
  0.006875,   0.006875,    0.006875,    0.006875,
  0.006875,   0.006875,    0.006875,    0.006875,
  0.006824,   0.006824,    0.006824,    0.006824,
  0.006803,   0.006803,    0.006803,    0.006803,
  0.006803,   0.006803,    0.006803,    0.006803,
  0.006792,   0.006792,    0.006792,    0.006792,
  0.006824,   0.006824,    0.006824,    0.006824,
  0.006835,   0.006835,    0.006835,    0.006835,
  0.006815,   0.006815,    0.006815,    0.006815,
  0.006795,   0.006795,    0.006795,    0.006795,
  0.006775,   0.006775,    0.006775,    0.006775,
  0.006755,   0.006755,    0.006755,    0.006755,
  0.006755,   0.006755,    0.006755,    0.006755,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006585,   0.006585,    0.006585,    0.006585,
  0.006385,   0.006385,    0.006385,    0.006385,
  0.006095,   0.006095,    0.006095,    0.006095,
  0.005819,   0.005819,    0.005819,    0.005819,
  0.00574,    0.00574,     0.00574,     0.00574,
  0.005663,   0.005663,    0.005663,    0.005663,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.00536,    0.00536,     0.00536,     0.00536,
  0.005377,   0.005377,    0.005377,    0.005377,
  0.00544,    0.00544,     0.00544,     0.00544,
  0.005525,   0.005525,    0.005525,    0.005525,
  0.005582,   0.005582,    0.005582,    0.005582,
  0.005551,   0.005551,    0.005551,    0.005551,
  0.005347,   0.005347,    0.005347,    0.005347,
  0.005032,   0.005032,    0.005032,    0.005032,
  0.004766,   0.004766,    0.004766,    0.004766,
  0.004611,   0.004611,    0.004611,    0.004611,
  0.004623,   0.004623,    0.004623,    0.004623,
  0.004675,   0.004675,    0.004675,    0.004675,
  0.004607,   0.004607,    0.004607,    0.004607,
  0.004577,   0.004577,    0.004577,    0.004577,
  0.004699,   0.004699,    0.004699,    0.004699,
  0.004748,   0.004748,    0.004748,    0.004748,
  0.004782,   0.004782,    0.004782,    0.004782,
  0.004786,   0.004786,    0.004786,    0.004786,
  0.004879,   0.004879,    0.004879,    0.004879,
  0.005108,   0.005108,    0.005108,    0.005108,
  0.005124,   0.005124,    0.005124,    0.005124,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.004857,   0.004857,    0.004857,    0.004857,
  0.0047,     0.0047,      0.0047,      0.0047,
  0.004544,   0.004544,    0.004544,    0.004544,
  0.004436,   0.004436,    0.004436,    0.004436,
  0.004391,   0.004391,    0.004391,    0.004391,
  0.004345,   0.004345,    0.004345,    0.004345,
  0.004267,   0.004267,    0.004267,    0.004267,
  0.004158,   0.004158,    0.004158,    0.004158,
  0.004046,   0.004046,    0.004046,    0.004046,
  0.003967,   0.003967,    0.003967,    0.003967,
  0.003918,   0.003918,    0.003918,    0.003918,
  0.003884,   0.003884,    0.003884,    0.003884,
  0.003897,   0.003897,    0.003897,    0.003897,
  0.003928,   0.003928,    0.003928,    0.003928,
  0.003911,   0.003911,    0.003911,    0.003911,
  0.003894,   0.003894,    0.003894,    0.003894,
  0.003878,   0.003878,    0.003878,    0.003878,
  0.003848,   0.003848,    0.003848,    0.003848,
  0.003884,   0.003884,    0.003884,    0.003884,
  0.003985,   0.003985,    0.003985,    0.003985,
  0.004055,   0.004055,    0.004055,    0.004055,
  0.004081,   0.004081,    0.004081,    0.004081,
  0.004122,   0.004122,    0.004122,    0.004122,
  0.004144,   0.004144,    0.004144,    0.004144,
  0.004152,   0.004152,    0.004152,    0.004152,
  0.004174,   0.004174,    0.004174,    0.004174,
  0.004178,   0.004178,    0.004178,    0.004178,
  0.004142,   0.004142,    0.004142,    0.004142,
  0.004121,   0.004121,    0.004121,    0.004121,
  0.004166,   0.004166,    0.004166,    0.004166,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004298,   0.004298,    0.004298,    0.004298,
  0.004342,   0.004342,    0.004342,    0.004342,
  0.004375,   0.004375,    0.004375,    0.004375,
  0.004384,   0.004384,    0.004384,    0.004384,
  0.004367,   0.004367,    0.004367,    0.004367,
  0.004293,   0.004293,    0.004293,    0.004293,
  0.004177,   0.004177,    0.004177,    0.004177,
  0.003944,   0.003944,    0.003944,    0.003944,
  0.003776,   0.003776,    0.003776,    0.003776,
  0.003701,   0.003701,    0.003701,    0.003701,
  0.003635,   0.003635,    0.003635,    0.003635,
  0.00354,    0.00354,     0.00354,     0.00354,
  0.00347,    0.00347,     0.00347,     0.00347,
  0.003436,   0.003436,    0.003436,    0.003436,
  0.003528,   0.003528,    0.003528,    0.003528,
  0.003724,   0.003724,    0.003724,    0.003724,
  0.003739,   0.003739,    0.003739,    0.003739,
  0.003747,   0.003747,    0.003747,    0.003747,
  0.003758,   0.003758,    0.003758,    0.003758,
  0.00378,    0.00378,     0.00378,     0.00378,
  0.00385,    0.00385,     0.00385,     0.00385,
  0.003851,   0.003851,    0.003851,    0.003851,
  0.003857,   0.003857,    0.003857,    0.003857,
  0.003839,   0.003839,    0.003839,    0.003839,
  0.00379,    0.00379,     0.00379,     0.00379,
  0.003872,   0.003872,    0.003872,    0.003872,
  0.003921,   0.003921,    0.003921,    0.003921,
  0.003853,   0.003853,    0.003853,    0.003853,
  0.003836,   0.003836,    0.003836,    0.003836,
  0.003848,   0.003848,    0.003848,    0.003848,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003984,   0.003984,    0.003984,    0.003984,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.004047,   0.004047,    0.004047,    0.004047,
  0.004073,   0.004073,    0.004073,    0.004073,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004567,   0.004567,    0.004567,    0.004567,
  0.004687,   0.004687,    0.004687,    0.004687,
  0.00462,    0.00462,     0.00462,     0.00462,
  0.00442,    0.00442,     0.00442,     0.00442,
  0.004257,   0.004257,    0.004257,    0.004257,
  0.004142,   0.004142,    0.004142,    0.004142,
  0.004019,   0.004019,    0.004019,    0.004019,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003936,   0.003936,    0.003936,    0.003936,
  0.004006,   0.004006,    0.004006,    0.004006,
  0.004041,   0.004041,    0.004041,    0.004041,
  0.004011,   0.004011,    0.004011,    0.004011,
  0.004115,   0.004115,    0.004115,    0.004115,
  0.004174,   0.004174,    0.004174,    0.004174,
  0.004205,   0.004205,    0.004205,    0.004205,
  0.004321,   0.004321,    0.004321,    0.004321,
  0.004384,   0.004384,    0.004384,    0.004384,
  0.004406,   0.004406,    0.004406,    0.004406,
  0.004409,   0.004409,    0.004409,    0.004409,
  0.004412,   0.004412,    0.004412,    0.004412,
  0.004405,   0.004405,    0.004405,    0.004405,
  0.004403,   0.004403,    0.004403,    0.004403,
  0.004423,   0.004423,    0.004423,    0.004423,
  0.004427,   0.004427,    0.004427,    0.004427,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.004473,   0.004473,    0.004473,    0.004473,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.00401,    0.00401,     0.00401,     0.00401,
  0.003922,   0.003922,    0.003922,    0.003922,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.003984,   0.003984,    0.003984,    0.003984,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004515,   0.004515,    0.004515,    0.004515,
  0.00464,    0.00464,     0.00464,     0.00464,
  0.004548,   0.004548,    0.004548,    0.004548,
  0.004352,   0.004352,    0.004352,    0.004352,
  0.00424,    0.00424,     0.00424,     0.00424,
  0.004162,   0.004162,    0.004162,    0.004162,
  0.004101,   0.004101,    0.004101,    0.004101,
  0.004025,   0.004025,    0.004025,    0.004025,
  0.003965,   0.003965,    0.003965,    0.003965,
  0.003933,   0.003933,    0.003933,    0.003933,
  0.00393,    0.00393,     0.00393,     0.00393,
  0.003944,   0.003944,    0.003944,    0.003944,
  0.003942,   0.003942,    0.003942,    0.003942,
  0.003894,   0.003894,    0.003894,    0.003894,
  0.003878,   0.003878,    0.003878,    0.003878,
  0.00388,    0.00388,     0.00388,     0.00388,
  0.003867,   0.003867,    0.003867,    0.003867,
  0.003869,   0.003869,    0.003869,    0.003869,
  0.003837,   0.003837,    0.003837,    0.003837,
  0.003839,   0.003839,    0.003839,    0.003839,
  0.003859,   0.003859,    0.003859,    0.003859,
  0.003881,   0.003881,    0.003881,    0.003881,
  0.003912,   0.003912,    0.003912,    0.003912,
  0.003828,   0.003828,    0.003828,    0.003828,
  0.003729,   0.003729,    0.003729,    0.003729,
  0.003761,   0.003761,    0.003761,    0.003761,
  0.003855,   0.003855,    0.003855,    0.003855,
  0.003902,   0.003902,    0.003902,    0.003902,
  0.003887,   0.003887,    0.003887,    0.003887,
  0.003887,   0.003887,    0.003887,    0.003887,
  0.004054,   0.004054,    0.004054,    0.004054,
  0.004226,   0.004226,    0.004226,    0.004226,
  0.004277,   0.004277,    0.004277,    0.004277,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004386,   0.004386,    0.004386,    0.004386,
  0.004361,   0.004361,    0.004361,    0.004361,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004333,   0.004333,    0.004333,    0.004333,
  0.004356,   0.004356,    0.004356,    0.004356,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004361,   0.004361,    0.004361,    0.004361,
  0.004424,   0.004424,    0.004424,    0.004424,
  0.004472,   0.004472,    0.004472,    0.004472,
  0.004487,   0.004487,    0.004487,    0.004487,
  0.004532,   0.004532,    0.004532,    0.004532,
  0.004623,   0.004623,    0.004623,    0.004623,
  0.004731,   0.004731,    0.004731,    0.004731,
  0.004855,   0.004855,    0.004855,    0.004855,
  0.004965,   0.004965,    0.004965,    0.004965,
  0.005076,   0.005076,    0.005076,    0.005076,
  0.005224,   0.005224,    0.005224,    0.005224,
  0.005342,   0.005342,    0.005342,    0.005342,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005441,   0.005441,    0.005441,    0.005441,
  0.005492,   0.005492,    0.005492,    0.005492,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.005484,   0.005484,    0.005484,    0.005484,
  0.005521,   0.005521,    0.005521,    0.005521,
  0.005559,   0.005559,    0.005559,    0.005559,
  0.005516,   0.005516,    0.005516,    0.005516,
  0.00544,    0.00544,     0.00544,     0.00544,
  0.005409,   0.005409,    0.005409,    0.005409,
  0.00539,    0.00539,     0.00539,     0.00539,
  0.005383,   0.005383,    0.005383,    0.005383,
  0.005389,   0.005389,    0.005389,    0.005389,
  0.005364,   0.005364,    0.005364,    0.005364,
  0.005326,   0.005326,    0.005326,    0.005326,
  0.005294,   0.005294,    0.005294,    0.005294,
  0.005231,   0.005231,    0.005231,    0.005231,
  0.005226,   0.005226,    0.005226,    0.005226,
  0.005257,   0.005257,    0.005257,    0.005257,
  0.00525,    0.00525,     0.00525,     0.00525,
  0.005244,   0.005244,    0.005244,    0.005244,
  0.005231,   0.005231,    0.005231,    0.005231,
  0.005269,   0.005269,    0.005269,    0.005269,
  0.005471,   0.005471,    0.005471,    0.005471,
  0.005762,   0.005762,    0.005762,    0.005762,
  0.005916,   0.005916,    0.005916,    0.005916,
  0.005974,   0.005974,    0.005974,    0.005974,
  0.006037,   0.006037,    0.006037,    0.006037,
  0.006105,   0.006105,    0.006105,    0.006105,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.006178,   0.006178,    0.006178,    0.006178,
  0.006234,   0.006234,    0.006234,    0.006234,
  0.006252,   0.006252,    0.006252,    0.006252,
  0.006252,   0.006252,    0.006252,    0.006252,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006384,   0.006384,    0.006384,    0.006384,
  0.006442,   0.006442,    0.006442,    0.006442,
  0.006507,   0.006507,    0.006507,    0.006507,
  0.006553,   0.006553,    0.006553,    0.006553,
  0.006604,   0.006604,    0.006604,    0.006604,
  0.006636,   0.006636,    0.006636,    0.006636,
  0.006672,   0.006672,    0.006672,    0.006672,
  0.006538,   0.006538,    0.006538,    0.006538,
  0.006199,   0.006199,    0.006199,    0.006199,
  0.005958,   0.005958,    0.005958,    0.005958,
  0.005958,   0.005958,    0.005958,    0.005958,
  0.005601,   0.005601,    0.005601,    0.005601,
  0.00488,    0.00488,     0.00488,     0.00488,
  0.004573,   0.004573,    0.004573,    0.004573,
  0.004498,   0.004498,    0.004498,    0.004498,
  0.004301,   0.004301,    0.004301,    0.004301,
  0.003986,   0.003986,    0.003986,    0.003986,
  0.003809,   0.003809,    0.003809,    0.003809,
  0.004079,   0.004079,    0.004079,    0.004079,
  0.004454,   0.004454,    0.004454,    0.004454,
  0.004403,   0.004403,    0.004403,    0.004403,
  0.004245,   0.004245,    0.004245,    0.004245,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.004146,   0.004146,    0.004146,    0.004146,
  0.004209,   0.004209,    0.004209,    0.004209,
  0.004304,   0.004304,    0.004304,    0.004304,
  0.004398,   0.004398,    0.004398,    0.004398,
  0.004382,   0.004382,    0.004382,    0.004382,
  0.004337,   0.004337,    0.004337,    0.004337,
  0.004291,   0.004291,    0.004291,    0.004291,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004225,   0.004225,    0.004225,    0.004225,
  0.004193,   0.004193,    0.004193,    0.004193,
  0.004177,   0.004177,    0.004177,    0.004177,
  0.00413,    0.00413,     0.00413,     0.00413,
  0.004067,   0.004067,    0.004067,    0.004067,
  0.004052,   0.004052,    0.004052,    0.004052,
  0.004052,   0.004052,    0.004052,    0.004052,
  0.004036,   0.004036,    0.004036,    0.004036,
  0.00402,    0.00402,     0.00402,     0.00402,
  0.004038,   0.004038,    0.004038,    0.004038,
  0.004071,   0.004071,    0.004071,    0.004071,
  0.004041,   0.004041,    0.004041,    0.004041,
  0.004026,   0.004026,    0.004026,    0.004026,
  0.004074,   0.004074,    0.004074,    0.004074,
  0.004063,   0.004063,    0.004063,    0.004063,
  0.00403,    0.00403,     0.00403,     0.00403,
  0.004018,   0.004018,    0.004018,    0.004018,
  0.003976,   0.003976,    0.003976,    0.003976,
  0.003945,   0.003945,    0.003945,    0.003945,
  0.003945,   0.003945,    0.003945,    0.003945,
  0.003944,   0.003944,    0.003944,    0.003944,
  0.004001,   0.004001,    0.004001,    0.004001,
  0.004088,   0.004088,    0.004088,    0.004088,
  0.004183,   0.004183,    0.004183,    0.004183,
  0.004209,   0.004209,    0.004209,    0.004209,
  0.004209,   0.004209,    0.004209,    0.004209,
  0.004244,   0.004244,    0.004244,    0.004244,
  0.004106,   0.004106,    0.004106,    0.004106,
  0.003918,   0.003918,    0.003918,    0.003918,
  0.003952,   0.003952,    0.003952,    0.003952,
  0.00408,    0.00408,     0.00408,     0.00408,
  0.004114,   0.004114,    0.004114,    0.004114,
  0.004131,   0.004131,    0.004131,    0.004131,
  0.004116,   0.004116,    0.004116,    0.004116,
  0.004087,   0.004087,    0.004087,    0.004087,
  0.004167,   0.004167,    0.004167,    0.004167,
  0.00423,    0.00423,     0.00423,     0.00423,
  0.004199,   0.004199,    0.004199,    0.004199,
  0.00409,    0.00409,     0.00409,     0.00409,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.004024,   0.004024,    0.004024,    0.004024,
  0.004056,   0.004056,    0.004056,    0.004056,
  0.004027,   0.004027,    0.004027,    0.004027,
  0.004016,   0.004016,    0.004016,    0.004016,
  0.004096,   0.004096,    0.004096,    0.004096,
  0.004212,   0.004212,    0.004212,    0.004212,
  0.004464,   0.004464,    0.004464,    0.004464,
  0.004912,   0.004912,    0.004912,    0.004912,
  0.005304,   0.005304,    0.005304,    0.005304,
  0.005563,   0.005563,    0.005563,    0.005563,
  0.005803,   0.005803,    0.005803,    0.005803,
  0.006009,   0.006009,    0.006009,    0.006009,
  0.005748,   0.005748,    0.005748,    0.005748,
  0.005332,   0.005332,    0.005332,    0.005332,
  0.005042,   0.005042,    0.005042,    0.005042,
  0.004773,   0.004773,    0.004773,    0.004773,
  0.004649,   0.004649,    0.004649,    0.004649,
  0.004408,   0.004408,    0.004408,    0.004408,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.003784,   0.003784,    0.003784,    0.003784,
  0.003624,   0.003624,    0.003624,    0.003624,
  0.003561,   0.003561,    0.003561,    0.003561,
  0.003498,   0.003498,    0.003498,    0.003498,
  0.003515,   0.003515,    0.003515,    0.003515,
  0.003564,   0.003564,    0.003564,    0.003564,
  0.003564,   0.003564,    0.003564,    0.003564,
  0.003515,   0.003515,    0.003515,    0.003515,
  0.003576,   0.003576,    0.003576,    0.003576,
  0.003687,   0.003687,    0.003687,    0.003687,
  0.003758,   0.003758,    0.003758,    0.003758,
  0.003865,   0.003865,    0.003865,    0.003865,
  0.004007,   0.004007,    0.004007,    0.004007,
  0.004057,   0.004057,    0.004057,    0.004057,
  0.004067,   0.004067,    0.004067,    0.004067,
  0.004148,   0.004148,    0.004148,    0.004148,
  0.004205,   0.004205,    0.004205,    0.004205,
  0.004306,   0.004306,    0.004306,    0.004306,
  0.004452,   0.004452,    0.004452,    0.004452,
  0.004585,   0.004585,    0.004585,    0.004585,
  0.004706,   0.004706,    0.004706,    0.004706,
  0.004734,   0.004734,    0.004734,    0.004734,
  0.004719,   0.004719,    0.004719,    0.004719,
  0.004725,   0.004725,    0.004725,    0.004725,
  0.004796,   0.004796,    0.004796,    0.004796,
  0.004945,   0.004945,    0.004945,    0.004945,
  0.005094,   0.005094,    0.005094,    0.005094,
  0.0052,     0.0052,      0.0052,      0.0052,
  0.005286,   0.005286,    0.005286,    0.005286,
  0.005349,   0.005349,    0.005349,    0.005349,
  0.00538,    0.00538,     0.00538,     0.00538,
  0.005372,   0.005372,    0.005372,    0.005372,
  0.005344,   0.005344,    0.005344,    0.005344,
  0.005336,   0.005336,    0.005336,    0.005336,
  0.005305,   0.005305,    0.005305,    0.005305,
  0.005242,   0.005242,    0.005242,    0.005242,
  0.005191,   0.005191,    0.005191,    0.005191,
  0.005183,   0.005183,    0.005183,    0.005183,
  0.005183,   0.005183,    0.005183,    0.005183,
  0.005215,   0.005215,    0.005215,    0.005215,
  0.005283,   0.005283,    0.005283,    0.005283,
  0.005327,   0.005327,    0.005327,    0.005327,
  0.005397,   0.005397,    0.005397,    0.005397,
  0.005479,   0.005479,    0.005479,    0.005479,
  0.00553,    0.00553,     0.00553,     0.00553,
  0.00553,    0.00553,     0.00553,     0.00553,
  0.005554,   0.005554,    0.005554,    0.005554,
  0.005617,   0.005617,    0.005617,    0.005617,
  0.005624,   0.005624,    0.005624,    0.005624,
  0.0056,     0.0056,      0.0056,      0.0056,
  0.005608,   0.005608,    0.005608,    0.005608,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005647,   0.005647,    0.005647,    0.005647,
  0.005699,   0.005699,    0.005699,    0.005699,
  0.00573,    0.00573,     0.00573,     0.00573,
  0.00575,    0.00575,     0.00575,     0.00575,
  0.00577,    0.00577,     0.00577,     0.00577,
  0.005758,   0.005758,    0.005758,    0.005758,
  0.005787,   0.005787,    0.005787,    0.005787,
  0.005816,   0.005816,    0.005816,    0.005816,
  0.005825,   0.005825,    0.005825,    0.005825,
  0.005897,   0.005897,    0.005897,    0.005897,
  0.00597,    0.00597,     0.00597,     0.00597,
  0.006132,   0.006132,    0.006132,    0.006132,
  0.00636,    0.00636,     0.00636,     0.00636,
  0.006478,   0.006478,    0.006478,    0.006478,
  0.006538,   0.006538,    0.006538,    0.006538,
  0.006563,   0.006563,    0.006563,    0.006563,
  0.006527,   0.006527,    0.006527,    0.006527,
  0.006483,   0.006483,    0.006483,    0.006483,
  0.006462,   0.006462,    0.006462,    0.006462,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.00641,    0.00641,     0.00641,     0.00641,
  0.006368,   0.006368,    0.006368,    0.006368,
  0.006326,   0.006326,    0.006326,    0.006326,
  0.006241,   0.006241,    0.006241,    0.006241,
  0.00618,    0.00618,     0.00618,     0.00618,
  0.006232,   0.006232,    0.006232,    0.006232,
  0.006325,   0.006325,    0.006325,    0.006325,
  0.006368,   0.006368,    0.006368,    0.006368,
  0.006368,   0.006368,    0.006368,    0.006368,
  0.006349,   0.006349,    0.006349,    0.006349,
  0.00631,    0.00631,     0.00631,     0.00631,
  0.006221,   0.006221,    0.006221,    0.006221,
  0.006176,   0.006176,    0.006176,    0.006176,
  0.00619,    0.00619,     0.00619,     0.00619,
  0.006128,   0.006128,    0.006128,    0.006128,
  0.006042,   0.006042,    0.006042,    0.006042,
  0.005969,   0.005969,    0.005969,    0.005969,
  0.005915,   0.005915,    0.005915,    0.005915,
  0.005875,   0.005875,    0.005875,    0.005875,
  0.005784,   0.005784,    0.005784,    0.005784,
  0.00568,    0.00568,     0.00568,     0.00568,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005614,   0.005614,    0.005614,    0.005614,
  0.005668,   0.005668,    0.005668,    0.005668,
  0.005706,   0.005706,    0.005706,    0.005706,
  0.005745,   0.005745,    0.005745,    0.005745,
  0.005834,   0.005834,    0.005834,    0.005834,
  0.005888,   0.005888,    0.005888,    0.005888,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005979,   0.005979,    0.005979,    0.005979,
  0.006021,   0.006021,    0.006021,    0.006021,
  0.006063,   0.006063,    0.006063,    0.006063,
  0.006157,   0.006157,    0.006157,    0.006157,
  0.006303,   0.006303,    0.006303,    0.006303,
  0.006451,   0.006451,    0.006451,    0.006451,
  0.006558,   0.006558,    0.006558,    0.006558,
  0.006665,   0.006665,    0.006665,    0.006665,
  0.006714,   0.006714,    0.006714,    0.006714,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006707,   0.006707,    0.006707,    0.006707,
  0.006658,   0.006658,    0.006658,    0.006658,
  0.006535,   0.006535,    0.006535,    0.006535,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.006419,   0.006419,    0.006419,    0.006419,
  0.006406,   0.006406,    0.006406,    0.006406,
  0.006404,   0.006404,    0.006404,    0.006404,
  0.00637,    0.00637,     0.00637,     0.00637,
  0.006316,   0.006316,    0.006316,    0.006316,
  0.006262,   0.006262,    0.006262,    0.006262,
  0.00623,    0.00623,     0.00623,     0.00623,
  0.006283,   0.006283,    0.006283,    0.006283,
  0.006367,   0.006367,    0.006367,    0.006367,
  0.006409,   0.006409,    0.006409,    0.006409,
  0.006335,   0.006335,    0.006335,    0.006335,
  0.006146,   0.006146,    0.006146,    0.006146,
  0.005957,   0.005957,    0.005957,    0.005957,
  0.005884,   0.005884,    0.005884,    0.005884,
  0.005947,   0.005947,    0.005947,    0.005947,
  0.00601,    0.00601,     0.00601,     0.00601,
  0.005989,   0.005989,    0.005989,    0.005989,
  0.005957,   0.005957,    0.005957,    0.005957,
  0.005926,   0.005926,    0.005926,    0.005926,
  0.005875,   0.005875,    0.005875,    0.005875,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.005724,   0.005724,    0.005724,    0.005724,
  0.005715,   0.005715,    0.005715,    0.005715,
  0.005711,   0.005711,    0.005711,    0.005711,
  0.005716,   0.005716,    0.005716,    0.005716,
  0.005704,   0.005704,    0.005704,    0.005704,
  0.005655,   0.005655,    0.005655,    0.005655,
  0.005609,   0.005609,    0.005609,    0.005609,
  0.005546,   0.005546,    0.005546,    0.005546,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.005475,   0.005475,    0.005475,    0.005475,
  0.005479,   0.005479,    0.005479,    0.005479,
  0.00551,    0.00551,     0.00551,     0.00551,
  0.005524,   0.005524,    0.005524,    0.005524,
  0.005548,   0.005548,    0.005548,    0.005548,
  0.005585,   0.005585,    0.005585,    0.005585,
  0.005629,   0.005629,    0.005629,    0.005629,
  0.005698,   0.005698,    0.005698,    0.005698,
  0.005747,   0.005747,    0.005747,    0.005747,
  0.005732,   0.005732,    0.005732,    0.005732,
  0.005612,   0.005612,    0.005612,    0.005612,
  0.005488,   0.005488,    0.005488,    0.005488,
  0.005439,   0.005439,    0.005439,    0.005439,
  0.00542,    0.00542,     0.00542,     0.00542,
  0.005342,   0.005342,    0.005342,    0.005342,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005319,   0.005319,    0.005319,    0.005319,
  0.005391,   0.005391,    0.005391,    0.005391,
  0.005431,   0.005431,    0.005431,    0.005431,
  0.005472,   0.005472,    0.005472,    0.005472,
  0.005481,   0.005481,    0.005481,    0.005481,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005638,   0.005638,    0.005638,    0.005638,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005738,   0.005738,    0.005738,    0.005738,
  0.005839,   0.005839,    0.005839,    0.005839,
  0.005929,   0.005929,    0.005929,    0.005929,
  0.005958,   0.005958,    0.005958,    0.005958,
  0.005936,   0.005936,    0.005936,    0.005936,
  0.005905,   0.005905,    0.005905,    0.005905,
  0.005884,   0.005884,    0.005884,    0.005884,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005821,   0.005821,    0.005821,    0.005821,
  0.00581,    0.00581,     0.00581,     0.00581,
  0.005821,   0.005821,    0.005821,    0.005821,
  0.005852,   0.005852,    0.005852,    0.005852,
  0.005863,   0.005863,    0.005863,    0.005863,
  0.005852,   0.005852,    0.005852,    0.005852,
  0.005831,   0.005831,    0.005831,    0.005831,
  0.005831,   0.005831,    0.005831,    0.005831,
  0.005842,   0.005842,    0.005842,    0.005842,
  0.005789,   0.005789,    0.005789,    0.005789,
  0.005726,   0.005726,    0.005726,    0.005726,
  0.005727,   0.005727,    0.005727,    0.005727,
  0.00577,    0.00577,     0.00577,     0.00577,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.005898,   0.005898,    0.005898,    0.005898,
  0.006244,   0.006244,    0.006244,    0.006244,
  0.006518,   0.006518,    0.006518,    0.006518,
  0.006538,   0.006538,    0.006538,    0.006538,
  0.006494,   0.006494,    0.006494,    0.006494,
  0.006546,   0.006546,    0.006546,    0.006546,
  0.006231,   0.006231,    0.006231,    0.006231,
  0.006016,   0.006016,    0.006016,    0.006016,
  0.006349,   0.006349,    0.006349,    0.006349,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.00575,    0.00575,     0.00575,     0.00575,
  0.005727,   0.005727,    0.005727,    0.005727,
  0.005806,   0.005806,    0.005806,    0.005806,
  0.005816,   0.005816,    0.005816,    0.005816,
  0.005699,   0.005699,    0.005699,    0.005699,
  0.005492,   0.005492,    0.005492,    0.005492,
  0.005175,   0.005175,    0.005175,    0.005175,
  0.005126,   0.005126,    0.005126,    0.005126,
  0.00544,    0.00544,     0.00544,     0.00544,
  0.005605,   0.005605,    0.005605,    0.005605,
  0.005659,   0.005659,    0.005659,    0.005659,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005401,   0.005401,    0.005401,    0.005401,
  0.005307,   0.005307,    0.005307,    0.005307,
  0.005263,   0.005263,    0.005263,    0.005263,
  0.005263,   0.005263,    0.005263,    0.005263,
  0.005332,   0.005332,    0.005332,    0.005332,
  0.005445,   0.005445,    0.005445,    0.005445,
  0.005439,   0.005439,    0.005439,    0.005439,
  0.005458,   0.005458,    0.005458,    0.005458,
  0.005718,   0.005718,    0.005718,    0.005718,
  0.006002,   0.006002,    0.006002,    0.006002,
  0.006202,   0.006202,    0.006202,    0.006202,
  0.006491,   0.006491,    0.006491,    0.006491,
  0.006803,   0.006803,    0.006803,    0.006803,
  0.006966,   0.006966,    0.006966,    0.006966,
  0.007072,   0.007072,    0.007072,    0.007072,
  0.00716,    0.00716,     0.00716,     0.00716,
  0.007179,   0.007179,    0.007179,    0.007179,
  0.0072,     0.0072,      0.0072,      0.0072,
  0.007295,   0.007295,    0.007295,    0.007295,
  0.007143,   0.007143,    0.007143,    0.007143,
  0.00665,    0.00665,     0.00665,     0.00665,
  0.006069,   0.006069,    0.006069,    0.006069,
  0.005622,   0.005622,    0.005622,    0.005622,
  0.005571,   0.005571,    0.005571,    0.005571,
  0.00568,    0.00568,     0.00568,     0.00568,
  0.005905,   0.005905,    0.005905,    0.005905,
  0.005981,   0.005981,    0.005981,    0.005981,
  0.005801,   0.005801,    0.005801,    0.005801,
  0.005753,   0.005753,    0.005753,    0.005753,
  0.005621,   0.005621,    0.005621,    0.005621,
  0.005582,   0.005582,    0.005582,    0.005582,
  0.005744,   0.005744,    0.005744,    0.005744,
  0.005758,   0.005758,    0.005758,    0.005758,
  0.005548,   0.005548,    0.005548,    0.005548,
  0.005437,   0.005437,    0.005437,    0.005437,
  0.005595,   0.005595,    0.005595,    0.005595,
  0.00574,    0.00574,     0.00574,     0.00574,
  0.005548,   0.005548,    0.005548,    0.005548,
  0.005305,   0.005305,    0.005305,    0.005305,
  0.005292,   0.005292,    0.005292,    0.005292,
  0.005382,   0.005382,    0.005382,    0.005382,
  0.005414,   0.005414,    0.005414,    0.005414,
  0.00536,    0.00536,     0.00536,     0.00536,
  0.00543,    0.00543,     0.00543,     0.00543,
  0.005449,   0.005449,    0.005449,    0.005449,
  0.005405,   0.005405,    0.005405,    0.005405,
  0.005394,   0.005394,    0.005394,    0.005394,
  0.005415,   0.005415,    0.005415,    0.005415,
  0.005468,   0.005468,    0.005468,    0.005468,
  0.00552,    0.00552,     0.00552,     0.00552,
  0.005539,   0.005539,    0.005539,    0.005539,
  0.005518,   0.005518,    0.005518,    0.005518,
  0.005454,   0.005454,    0.005454,    0.005454,
  0.00538,    0.00538,     0.00538,     0.00538,
  0.005402,   0.005402,    0.005402,    0.005402,
  0.005486,   0.005486,    0.005486,    0.005486,
  0.005633,   0.005633,    0.005633,    0.005633,
  0.005759,   0.005759,    0.005759,    0.005759,
  0.006037,   0.006037,    0.006037,    0.006037,
  0.006341,   0.006341,    0.006341,    0.006341,
  0.006274,   0.006274,    0.006274,    0.006274,
  0.006158,   0.006158,    0.006158,    0.006158,
  0.006195,   0.006195,    0.006195,    0.006195,
  0.00624,    0.00624,     0.00624,     0.00624,
  0.006286,   0.006286,    0.006286,    0.006286,
  0.00623,    0.00623,     0.00623,     0.00623,
  0.006132,   0.006132,    0.006132,    0.006132,
  0.006045,   0.006045,    0.006045,    0.006045,
  0.005931,   0.005931,    0.005931,    0.005931,
  0.00586,    0.00586,     0.00586,     0.00586,
  0.005807,   0.005807,    0.005807,    0.005807,
  0.005647,   0.005647,    0.005647,    0.005647,
  0.005364,   0.005364,    0.005364,    0.005364,
  0.005165,   0.005165,    0.005165,    0.005165,
  0.005083,   0.005083,    0.005083,    0.005083,
  0.005021,   0.005021,    0.005021,    0.005021,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.005031,   0.005031,    0.005031,    0.005031,
  0.005056,   0.005056,    0.005056,    0.005056,
  0.005119,   0.005119,    0.005119,    0.005119,
  0.005183,   0.005183,    0.005183,    0.005183,
  0.005034,   0.005034,    0.005034,    0.005034,
  0.00491,    0.00491,     0.00491,     0.00491,
  0.004933,   0.004933,    0.004933,    0.004933,
  0.004989,   0.004989,    0.004989,    0.004989,
  0.005234,   0.005234,    0.005234,    0.005234,
  0.005311,   0.005311,    0.005311,    0.005311,
  0.005191,   0.005191,    0.005191,    0.005191,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005445,   0.005445,    0.005445,    0.005445,
  0.005421,   0.005421,    0.005421,    0.005421,
  0.005182,   0.005182,    0.005182,    0.005182,
  0.005088,   0.005088,    0.005088,    0.005088,
  0.005089,   0.005089,    0.005089,    0.005089,
  0.005064,   0.005064,    0.005064,    0.005064,
  0.005036,   0.005036,    0.005036,    0.005036,
  0.005016,   0.005016,    0.005016,    0.005016,
  0.005081,   0.005081,    0.005081,    0.005081,
  0.005161,   0.005161,    0.005161,    0.005161,
  0.005221,   0.005221,    0.005221,    0.005221,
  0.005259,   0.005259,    0.005259,    0.005259,
  0.005248,   0.005248,    0.005248,    0.005248,
  0.005288,   0.005288,    0.005288,    0.005288,
  0.005324,   0.005324,    0.005324,    0.005324,
  0.00527,    0.00527,     0.00527,     0.00527,
  0.005252,   0.005252,    0.005252,    0.005252,
  0.005285,   0.005285,    0.005285,    0.005285,
  0.005351,   0.005351,    0.005351,    0.005351,
  0.005416,   0.005416,    0.005416,    0.005416,
  0.005416,   0.005416,    0.005416,    0.005416,
  0.005384,   0.005384,    0.005384,    0.005384,
  0.005336,   0.005336,    0.005336,    0.005336,
  0.005288,   0.005288,    0.005288,    0.005288,
  0.005256,   0.005256,    0.005256,    0.005256,
  0.00516,    0.00516,     0.00516,     0.00516,
  0.005015,   0.005015,    0.005015,    0.005015,
  0.004902,   0.004902,    0.004902,    0.004902,
  0.00473,    0.00473,     0.00473,     0.00473,
  0.004562,   0.004562,    0.004562,    0.004562,
  0.004509,   0.004509,    0.004509,    0.004509,
  0.004496,   0.004496,    0.004496,    0.004496,
  0.004513,   0.004513,    0.004513,    0.004513,
  0.004473,   0.004473,    0.004473,    0.004473,
  0.004402,   0.004402,    0.004402,    0.004402,
  0.004378,   0.004378,    0.004378,    0.004378,
  0.004368,   0.004368,    0.004368,    0.004368,
  0.004368,   0.004368,    0.004368,    0.004368,
  0.004406,   0.004406,    0.004406,    0.004406,
  0.004544,   0.004544,    0.004544,    0.004544,
  0.004701,   0.004701,    0.004701,    0.004701,
  0.004728,   0.004728,    0.004728,    0.004728,
  0.004791,   0.004791,    0.004791,    0.004791,
  0.004935,   0.004935,    0.004935,    0.004935,
  0.005022,   0.005022,    0.005022,    0.005022,
  0.005022,   0.005022,    0.005022,    0.005022,
  0.005038,   0.005038,    0.005038,    0.005038,
  0.005024,   0.005024,    0.005024,    0.005024,
  0.004818,   0.004818,    0.004818,    0.004818,
  0.004564,   0.004564,    0.004564,    0.004564,
  0.004494,   0.004494,    0.004494,    0.004494,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.004463,   0.004463,    0.004463,    0.004463,
  0.004444,   0.004444,    0.004444,    0.004444,
  0.004489,   0.004489,    0.004489,    0.004489,
  0.004616,   0.004616,    0.004616,    0.004616,
  0.004669,   0.004669,    0.004669,    0.004669,
  0.004655,   0.004655,    0.004655,    0.004655,
  0.004646,   0.004646,    0.004646,    0.004646,
  0.004534,   0.004534,    0.004534,    0.004534,
  0.004408,   0.004408,    0.004408,    0.004408,
  0.004373,   0.004373,    0.004373,    0.004373,
  0.004432,   0.004432,    0.004432,    0.004432,
  0.004513,   0.004513,    0.004513,    0.004513,
  0.004493,   0.004493,    0.004493,    0.004493,
  0.00448,    0.00448,     0.00448,     0.00448,
  0.004548,   0.004548,    0.004548,    0.004548,
  0.004588,   0.004588,    0.004588,    0.004588,
  0.004547,   0.004547,    0.004547,    0.004547,
  0.004511,   0.004511,    0.004511,    0.004511,
  0.004511,   0.004511,    0.004511,    0.004511,
  0.004475,   0.004475,    0.004475,    0.004475,
  0.004485,   0.004485,    0.004485,    0.004485,
  0.004544,   0.004544,    0.004544,    0.004544,
  0.00459,    0.00459,     0.00459,     0.00459,
  0.004639,   0.004639,    0.004639,    0.004639,
  0.004656,   0.004656,    0.004656,    0.004656,
  0.004639,   0.004639,    0.004639,    0.004639,
  0.004635,   0.004635,    0.004635,    0.004635,
  0.004663,   0.004663,    0.004663,    0.004663,
  0.00466,    0.00466,     0.00466,     0.00466,
  0.004657,   0.004657,    0.004657,    0.004657,
  0.00464,    0.00464,     0.00464,     0.00464,
  0.004591,   0.004591,    0.004591,    0.004591,
  0.004543,   0.004543,    0.004543,    0.004543,
  0.004497,   0.004497,    0.004497,    0.004497,
  0.004457,   0.004457,    0.004457,    0.004457,
  0.004368,   0.004368,    0.004368,    0.004368,
  0.004232,   0.004232,    0.004232,    0.004232,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004058,   0.004058,    0.004058,    0.004058,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003976,   0.003976,    0.003976,    0.003976,
  0.003977,   0.003977,    0.003977,    0.003977,
  0.003849,   0.003849,    0.003849,    0.003849,
  0.003719,   0.003719,    0.003719,    0.003719,
  0.00354,    0.00354,     0.00354,     0.00354,
  0.003456,   0.003456,    0.003456,    0.003456,
  0.003382,   0.003382,    0.003382,    0.003382,
  0.00304,    0.00304,     0.00304,     0.00304,
  0.002913,   0.002913,    0.002913,    0.002913,
  0.003058,   0.003058,    0.003058,    0.003058,
  0.002951,   0.002951,    0.002951,    0.002951,
  0.002732,   0.002732,    0.002732,    0.002732,
  0.002686,   0.002686,    0.002686,    0.002686,
  0.002823,   0.002823,    0.002823,    0.002823,
  0.003037,   0.003037,    0.003037,    0.003037,
  0.003182,   0.003182,    0.003182,    0.003182,
  0.003334,   0.003334,    0.003334,    0.003334,
  0.003528,   0.003528,    0.003528,    0.003528,
  0.003691,   0.003691,    0.003691,    0.003691,
  0.003927,   0.003927,    0.003927,    0.003927,
  0.00428,    0.00428,     0.00428,     0.00428,
  0.004676,   0.004676,    0.004676,    0.004676,
  0.005066,   0.005066,    0.005066,    0.005066,
  0.00547,    0.00547,     0.00547,     0.00547,
  0.005956,   0.005956,    0.005956,    0.005956,
  0.006354,   0.006354,    0.006354,    0.006354,
  0.006499,   0.006499,    0.006499,    0.006499,
  0.006518,   0.006518,    0.006518,    0.006518,
  0.006518,   0.006518,    0.006518,    0.006518,
  0.006518,   0.006518,    0.006518,    0.006518,
  0.006468,   0.006468,    0.006468,    0.006468,
  0.006328,   0.006328,    0.006328,    0.006328,
  0.006146,   0.006146,    0.006146,    0.006146,
  0.005974,   0.005974,    0.005974,    0.005974,
  0.005791,   0.005791,    0.005791,    0.005791,
  0.005583,   0.005583,    0.005583,    0.005583,
  0.005429,   0.005429,    0.005429,    0.005429,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005186,   0.005186,    0.005186,    0.005186,
  0.005379,   0.005379,    0.005379,    0.005379,
  0.005553,   0.005553,    0.005553,    0.005553,
  0.005602,   0.005602,    0.005602,    0.005602,
  0.005523,   0.005523,    0.005523,    0.005523,
  0.005334,   0.005334,    0.005334,    0.005334,
  0.005152,   0.005152,    0.005152,    0.005152,
  0.005097,   0.005097,    0.005097,    0.005097,
  0.00511,    0.00511,     0.00511,     0.00511,
  0.004939,   0.004939,    0.004939,    0.004939,
  0.004599,   0.004599,    0.004599,    0.004599,
  0.004523,   0.004523,    0.004523,    0.004523,
  0.004565,   0.004565,    0.004565,    0.004565,
  0.004343,   0.004343,    0.004343,    0.004343,
  0.004381,   0.004381,    0.004381,    0.004381,
  0.00491,    0.00491,     0.00491,     0.00491,
  0.005212,   0.005212,    0.005212,    0.005212,
  0.005184,   0.005184,    0.005184,    0.005184,
  0.005175,   0.005175,    0.005175,    0.005175,
  0.005266,   0.005266,    0.005266,    0.005266,
  0.005423,   0.005423,    0.005423,    0.005423,
  0.005581,   0.005581,    0.005581,    0.005581,
  0.005675,   0.005675,    0.005675,    0.005675,
  0.00572,    0.00572,     0.00572,     0.00572,
  0.005778,   0.005778,    0.005778,    0.005778,
  0.005931,   0.005931,    0.005931,    0.005931,
  0.006063,   0.006063,    0.006063,    0.006063,
  0.006126,   0.006126,    0.006126,    0.006126,
  0.006269,   0.006269,    0.006269,    0.006269,
  0.006404,   0.006404,    0.006404,    0.006404,
  0.006413,   0.006413,    0.006413,    0.006413,
  0.006399,   0.006399,    0.006399,    0.006399,
  0.00643,    0.00643,     0.00643,     0.00643,
  0.006462,   0.006462,    0.006462,    0.006462,
  0.006471,   0.006471,    0.006471,    0.006471,
  0.006439,   0.006439,    0.006439,    0.006439,
  0.006385,   0.006385,    0.006385,    0.006385,
  0.006354,   0.006354,    0.006354,    0.006354,
  0.006295,   0.006295,    0.006295,    0.006295,
  0.006255,   0.006255,    0.006255,    0.006255,
  0.006273,   0.006273,    0.006273,    0.006273,
  0.006291,   0.006291,    0.006291,    0.006291,
  0.006287,   0.006287,    0.006287,    0.006287,
  0.006324,   0.006324,    0.006324,    0.006324,
  0.006394,   0.006394,    0.006394,    0.006394,
  0.006413,   0.006413,    0.006413,    0.006413,
  0.006413,   0.006413,    0.006413,    0.006413,
  0.006445,   0.006445,    0.006445,    0.006445,
  0.006508,   0.006508,    0.006508,    0.006508,
  0.00653,    0.00653,     0.00653,     0.00653,
  0.00651,    0.00651,     0.00651,     0.00651,
  0.00646,    0.00646,     0.00646,     0.00646,
  0.006378,   0.006378,    0.006378,    0.006378,
  0.006314,   0.006314,    0.006314,    0.006314,
  0.006258,   0.006258,    0.006258,    0.006258,
  0.006225,   0.006225,    0.006225,    0.006225,
  0.006281,   0.006281,    0.006281,    0.006281,
  0.006499,   0.006499,    0.006499,    0.006499,
  0.00681,    0.00681,     0.00681,     0.00681,
  0.007034,   0.007034,    0.007034,    0.007034,
  0.007109,   0.007109,    0.007109,    0.007109,
  0.007182,   0.007182,    0.007182,    0.007182,
  0.00699,    0.00699,     0.00699,     0.00699,
  0.006374,   0.006374,    0.006374,    0.006374,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.005565,   0.005565,    0.005565,    0.005565,
  0.005502,   0.005502,    0.005502,    0.005502,
  0.005431,   0.005431,    0.005431,    0.005431,
  0.005384,   0.005384,    0.005384,    0.005384,
  0.00536,    0.00536,     0.00536,     0.00536,
  0.005344,   0.005344,    0.005344,    0.005344,
  0.005289,   0.005289,    0.005289,    0.005289,
  0.005245,   0.005245,    0.005245,    0.005245,
  0.005202,   0.005202,    0.005202,    0.005202,
  0.005196,   0.005196,    0.005196,    0.005196,
  0.005248,   0.005248,    0.005248,    0.005248,
  0.005286,   0.005286,    0.005286,    0.005286,
  0.005251,   0.005251,    0.005251,    0.005251,
  0.00523,    0.00523,     0.00523,     0.00523,
  0.005227,   0.005227,    0.005227,    0.005227,
  0.005161,   0.005161,    0.005161,    0.005161,
  0.005049,   0.005049,    0.005049,    0.005049,
  0.004938,   0.004938,    0.004938,    0.004938,
  0.004809,   0.004809,    0.004809,    0.004809,
  0.004649,   0.004649,    0.004649,    0.004649,
  0.004534,   0.004534,    0.004534,    0.004534,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004477,   0.004477,    0.004477,    0.004477,
  0.004366,   0.004366,    0.004366,    0.004366,
  0.004288,   0.004288,    0.004288,    0.004288,
  0.004195,   0.004195,    0.004195,    0.004195,
  0.004135,   0.004135,    0.004135,    0.004135,
  0.004137,   0.004137,    0.004137,    0.004137,
  0.004169,   0.004169,    0.004169,    0.004169,
  0.004185,   0.004185,    0.004185,    0.004185,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004214,   0.004214,    0.004214,    0.004214,
  0.004274,   0.004274,    0.004274,    0.004274,
  0.004354,   0.004354,    0.004354,    0.004354,
  0.004396,   0.004396,    0.004396,    0.004396,
  0.004434,   0.004434,    0.004434,    0.004434,
  0.004386,   0.004386,    0.004386,    0.004386,
  0.004186,   0.004186,    0.004186,    0.004186,
  0.003956,   0.003956,    0.003956,    0.003956,
  0.003766,   0.003766,    0.003766,    0.003766,
  0.003569,   0.003569,    0.003569,    0.003569,
  0.003355,   0.003355,    0.003355,    0.003355,
  0.003208,   0.003208,    0.003208,    0.003208,
  0.003175,   0.003175,    0.003175,    0.003175,
  0.003271,   0.003271,    0.003271,    0.003271,
  0.003357,   0.003357,    0.003357,    0.003357,
  0.003422,   0.003422,    0.003422,    0.003422,
  0.003582,   0.003582,    0.003582,    0.003582,
  0.003734,   0.003734,    0.003734,    0.003734,
  0.003805,   0.003805,    0.003805,    0.003805,
  0.003808,   0.003808,    0.003808,    0.003808,
  0.003738,   0.003738,    0.003738,    0.003738,
  0.003601,   0.003601,    0.003601,    0.003601,
  0.003549,   0.003549,    0.003549,    0.003549,
  0.003607,   0.003607,    0.003607,    0.003607,
  0.003768,   0.003768,    0.003768,    0.003768,
  0.003916,   0.003916,    0.003916,    0.003916,
  0.004049,   0.004049,    0.004049,    0.004049,
  0.004166,   0.004166,    0.004166,    0.004166,
  0.004165,   0.004165,    0.004165,    0.004165,
  0.00418,    0.00418,     0.00418,     0.00418,
  0.004257,   0.004257,    0.004257,    0.004257,
  0.00432,    0.00432,     0.00432,     0.00432,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004366,   0.004366,    0.004366,    0.004366,
  0.004429,   0.004429,    0.004429,    0.004429,
  0.004461,   0.004461,    0.004461,    0.004461,
  0.00443,    0.00443,     0.00443,     0.00443,
  0.004367,   0.004367,    0.004367,    0.004367,
  0.004273,   0.004273,    0.004273,    0.004273,
  0.004212,   0.004212,    0.004212,    0.004212,
  0.004217,   0.004217,    0.004217,    0.004217,
  0.00424,    0.00424,     0.00424,     0.00424,
  0.004216,   0.004216,    0.004216,    0.004216,
  0.004224,   0.004224,    0.004224,    0.004224,
  0.004266,   0.004266,    0.004266,    0.004266,
  0.00427,    0.00427,     0.00427,     0.00427,
  0.004252,   0.004252,    0.004252,    0.004252,
  0.004259,   0.004259,    0.004259,    0.004259,
  0.004366,   0.004366,    0.004366,    0.004366,
  0.004482,   0.004482,    0.004482,    0.004482,
  0.004545,   0.004545,    0.004545,    0.004545,
  0.004607,   0.004607,    0.004607,    0.004607,
  0.004704,   0.004704,    0.004704,    0.004704,
  0.004836,   0.004836,    0.004836,    0.004836,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.005157,   0.005157,    0.005157,    0.005157,
  0.005267,   0.005267,    0.005267,    0.005267,
  0.005307,   0.005307,    0.005307,    0.005307,
  0.005328,   0.005328,    0.005328,    0.005328,
  0.005372,   0.005372,    0.005372,    0.005372,
  0.005449,   0.005449,    0.005449,    0.005449,
  0.005556,   0.005556,    0.005556,    0.005556,
  0.005685,   0.005685,    0.005685,    0.005685,
  0.00581,    0.00581,     0.00581,     0.00581,
  0.005864,   0.005864,    0.005864,    0.005864,
  0.005922,   0.005922,    0.005922,    0.005922,
  0.005981,   0.005981,    0.005981,    0.005981,
  0.006016,   0.006016,    0.006016,    0.006016,
  0.006107,   0.006107,    0.006107,    0.006107,
  0.006168,   0.006168,    0.006168,    0.006168,
  0.006199,   0.006199,    0.006199,    0.006199,
  0.006241,   0.006241,    0.006241,    0.006241,
  0.006294,   0.006294,    0.006294,    0.006294,
  0.006336,   0.006336,    0.006336,    0.006336,
  0.006337,   0.006337,    0.006337,    0.006337,
  0.006338,   0.006338,    0.006338,    0.006338,
  0.00634,    0.00634,     0.00634,     0.00634,
  0.006334,   0.006334,    0.006334,    0.006334,
  0.006348,   0.006348,    0.006348,    0.006348,
  0.006384,   0.006384,    0.006384,    0.006384,
  0.006407,   0.006407,    0.006407,    0.006407,
  0.006381,   0.006381,    0.006381,    0.006381,
  0.006297,   0.006297,    0.006297,    0.006297,
  0.006214,   0.006214,    0.006214,    0.006214,
  0.006202,   0.006202,    0.006202,    0.006202,
  0.006178,   0.006178,    0.006178,    0.006178,
  0.006105,   0.006105,    0.006105,    0.006105,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006086,   0.006086,    0.006086,    0.006086,
  0.006123,   0.006123,    0.006123,    0.006123,
  0.006197,   0.006197,    0.006197,    0.006197,
  0.006328,   0.006328,    0.006328,    0.006328,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.006605,   0.006605,    0.006605,    0.006605,
  0.006692,   0.006692,    0.006692,    0.006692,
  0.00677,    0.00677,     0.00677,     0.00677,
  0.006777,   0.006777,    0.006777,    0.006777,
  0.006609,   0.006609,    0.006609,    0.006609,
  0.006517,   0.006517,    0.006517,    0.006517,
  0.006548,   0.006548,    0.006548,    0.006548,
  0.00643,    0.00643,     0.00643,     0.00643,
  0.006283,   0.006283,    0.006283,    0.006283,
  0.006073,   0.006073,    0.006073,    0.006073,
  0.005821,   0.005821,    0.005821,    0.005821,
  0.005634,   0.005634,    0.005634,    0.005634,
  0.00549,    0.00549,     0.00549,     0.00549,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005333,   0.005333,    0.005333,    0.005333,
  0.005311,   0.005311,    0.005311,    0.005311,
  0.005319,   0.005319,    0.005319,    0.005319,
  0.00536,    0.00536,     0.00536,     0.00536,
  0.005414,   0.005414,    0.005414,    0.005414,
  0.005468,   0.005468,    0.005468,    0.005468,
  0.005511,   0.005511,    0.005511,    0.005511,
  0.005605,   0.005605,    0.005605,    0.005605,
  0.005703,   0.005703,    0.005703,    0.005703,
  0.005785,   0.005785,    0.005785,    0.005785,
  0.005789,   0.005789,    0.005789,    0.005789,
  0.005743,   0.005743,    0.005743,    0.005743,
  0.005736,   0.005736,    0.005736,    0.005736,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005403,   0.005403,    0.005403,    0.005403,
  0.005353,   0.005353,    0.005353,    0.005353,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005296,   0.005296,    0.005296,    0.005296,
  0.005242,   0.005242,    0.005242,    0.005242,
  0.005188,   0.005188,    0.005188,    0.005188,
  0.005164,   0.005164,    0.005164,    0.005164,
  0.005204,   0.005204,    0.005204,    0.005204,
  0.005258,   0.005258,    0.005258,    0.005258,
  0.005321,   0.005321,    0.005321,    0.005321,
  0.005466,   0.005466,    0.005466,    0.005466,
  0.005623,   0.005623,    0.005623,    0.005623,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005697,   0.005697,    0.005697,    0.005697,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005766,   0.005766,    0.005766,    0.005766,
  0.005818,   0.005818,    0.005818,    0.005818,
  0.005836,   0.005836,    0.005836,    0.005836,
  0.005801,   0.005801,    0.005801,    0.005801,
  0.005748,   0.005748,    0.005748,    0.005748,
  0.005714,   0.005714,    0.005714,    0.005714,
  0.005724,   0.005724,    0.005724,    0.005724,
  0.005736,   0.005736,    0.005736,    0.005736,
  0.005604,   0.005604,    0.005604,    0.005604,
  0.005423,   0.005423,    0.005423,    0.005423,
  0.005295,   0.005295,    0.005295,    0.005295,
  0.005077,   0.005077,    0.005077,    0.005077,
  0.004866,   0.004866,    0.004866,    0.004866,
  0.00475,    0.00475,     0.00475,     0.00475,
  0.004687,   0.004687,    0.004687,    0.004687,
  0.004635,   0.004635,    0.004635,    0.004635,
  0.004593,   0.004593,    0.004593,    0.004593,
  0.004604,   0.004604,    0.004604,    0.004604,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004541,   0.004541,    0.004541,    0.004541,
  0.004491,   0.004491,    0.004491,    0.004491,
  0.004387,   0.004387,    0.004387,    0.004387,
  0.004362,   0.004362,    0.004362,    0.004362,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004426,   0.004426,    0.004426,    0.004426,
  0.004436,   0.004436,    0.004436,    0.004436,
  0.004426,   0.004426,    0.004426,    0.004426,
  0.004428,   0.004428,    0.004428,    0.004428,
  0.004419,   0.004419,    0.004419,    0.004419,
  0.004385,   0.004385,    0.004385,    0.004385,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004287,   0.004287,    0.004287,    0.004287,
  0.004272,   0.004272,    0.004272,    0.004272,
  0.004351,   0.004351,    0.004351,    0.004351,
  0.00443,    0.00443,     0.00443,     0.00443,
  0.004479,   0.004479,    0.004479,    0.004479,
  0.004606,   0.004606,    0.004606,    0.004606,
  0.004717,   0.004717,    0.004717,    0.004717,
  0.004764,   0.004764,    0.004764,    0.004764,
  0.004782,   0.004782,    0.004782,    0.004782,
  0.004815,   0.004815,    0.004815,    0.004815,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004714,   0.004714,    0.004714,    0.004714,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.005613,   0.005613,    0.005613,    0.005613,
  0.005806,   0.005806,    0.005806,    0.005806,
  0.0059,     0.0059,      0.0059,      0.0059,
  0.006011,   0.006011,    0.006011,    0.006011,
  0.006111,   0.006111,    0.006111,    0.006111,
  0.006128,   0.006128,    0.006128,    0.006128,
  0.006039,   0.006039,    0.006039,    0.006039,
  0.005864,   0.005864,    0.005864,    0.005864,
  0.005746,   0.005746,    0.005746,    0.005746,
  0.005727,   0.005727,    0.005727,    0.005727,
  0.005737,   0.005737,    0.005737,    0.005737,
  0.005737,   0.005737,    0.005737,    0.005737,
  0.005686,   0.005686,    0.005686,    0.005686,
  0.005585,   0.005585,    0.005585,    0.005585,
  0.005397,   0.005397,    0.005397,    0.005397,
  0.005327,   0.005327,    0.005327,    0.005327,
  0.005402,   0.005402,    0.005402,    0.005402,
  0.005468,   0.005468,    0.005468,    0.005468,
  0.005526,   0.005526,    0.005526,    0.005526,
  0.005531,   0.005531,    0.005531,    0.005531,
  0.005534,   0.005534,    0.005534,    0.005534,
  0.005518,   0.005518,    0.005518,    0.005518,
  0.005504,   0.005504,    0.005504,    0.005504,
  0.005465,   0.005465,    0.005465,    0.005465,
  0.005413,   0.005413,    0.005413,    0.005413,
  0.005335,   0.005335,    0.005335,    0.005335,
  0.005238,   0.005238,    0.005238,    0.005238,
  0.005215,   0.005215,    0.005215,    0.005215,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005131,   0.005131,    0.005131,    0.005131,
  0.005143,   0.005143,    0.005143,    0.005143,
  0.005137,   0.005137,    0.005137,    0.005137,
  0.005162,   0.005162,    0.005162,    0.005162,
  0.0052,     0.0052,      0.0052,      0.0052,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005259,   0.005259,    0.005259,    0.005259,
  0.005272,   0.005272,    0.005272,    0.005272,
  0.005299,   0.005299,    0.005299,    0.005299,
  0.005303,   0.005303,    0.005303,    0.005303,
  0.005318,   0.005318,    0.005318,    0.005318,
  0.005307,   0.005307,    0.005307,    0.005307,
  0.005284,   0.005284,    0.005284,    0.005284,
  0.005279,   0.005279,    0.005279,    0.005279,
  0.005262,   0.005262,    0.005262,    0.005262,
  0.005244,   0.005244,    0.005244,    0.005244,
  0.005241,   0.005241,    0.005241,    0.005241,
  0.005277,   0.005277,    0.005277,    0.005277,
  0.005365,   0.005365,    0.005365,    0.005365,
  0.005463,   0.005463,    0.005463,    0.005463,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005675,   0.005675,    0.005675,    0.005675,
  0.005788,   0.005788,    0.005788,    0.005788,
  0.005843,   0.005843,    0.005843,    0.005843,
  0.005962,   0.005962,    0.005962,    0.005962,
  0.006099,   0.006099,    0.006099,    0.006099,
  0.006215,   0.006215,    0.006215,    0.006215,
  0.00626,    0.00626,     0.00626,     0.00626,
  0.006211,   0.006211,    0.006211,    0.006211,
  0.006208,   0.006208,    0.006208,    0.006208,
  0.006273,   0.006273,    0.006273,    0.006273,
  0.006321,   0.006321,    0.006321,    0.006321,
  0.006312,   0.006312,    0.006312,    0.006312,
  0.006288,   0.006288,    0.006288,    0.006288,
  0.006248,   0.006248,    0.006248,    0.006248,
  0.006178,   0.006178,    0.006178,    0.006178,
  0.006175,   0.006175,    0.006175,    0.006175,
  0.006212,   0.006212,    0.006212,    0.006212,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.006095,   0.006095,    0.006095,    0.006095,
  0.005985,   0.005985,    0.005985,    0.005985,
  0.00588,    0.00588,     0.00588,     0.00588,
  0.005863,   0.005863,    0.005863,    0.005863,
  0.005868,   0.005868,    0.005868,    0.005868,
  0.005869,   0.005869,    0.005869,    0.005869,
  0.005858,   0.005858,    0.005858,    0.005858,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.005926,   0.005926,    0.005926,    0.005926,
  0.005898,   0.005898,    0.005898,    0.005898,
  0.005901,   0.005901,    0.005901,    0.005901,
  0.005897,   0.005897,    0.005897,    0.005897,
  0.00591,    0.00591,     0.00591,     0.00591,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.005906,   0.005906,    0.005906,    0.005906,
  0.005871,   0.005871,    0.005871,    0.005871,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005836,   0.005836,    0.005836,    0.005836,
  0.005801,   0.005801,    0.005801,    0.005801,
  0.005748,   0.005748,    0.005748,    0.005748,
  0.00568,    0.00568,     0.00568,     0.00568,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.006035,   0.006035,    0.006035,    0.006035,
  0.00608,    0.00608,     0.00608,     0.00608,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.006059,   0.006059,    0.006059,    0.006059,
  0.005973,   0.005973,    0.005973,    0.005973,
  0.005792,   0.005792,    0.005792,    0.005792,
  0.005721,   0.005721,    0.005721,    0.005721,
  0.005755,   0.005755,    0.005755,    0.005755,
  0.005671,   0.005671,    0.005671,    0.005671,
  0.005531,   0.005531,    0.005531,    0.005531,
  0.005499,   0.005499,    0.005499,    0.005499,
  0.005433,   0.005433,    0.005433,    0.005433,
  0.00539,    0.00539,     0.00539,     0.00539,
  0.005424,   0.005424,    0.005424,    0.005424,
  0.005448,   0.005448,    0.005448,    0.005448,
  0.00555,    0.00555,     0.00555,     0.00555,
  0.005729,   0.005729,    0.005729,    0.005729,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005935,   0.005935,    0.005935,    0.005935,
  0.006015,   0.006015,    0.006015,    0.006015,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.006013,   0.006013,    0.006013,    0.006013,
  0.005963,   0.005963,    0.005963,    0.005963,
  0.005894,   0.005894,    0.005894,    0.005894,
  0.005826,   0.005826,    0.005826,    0.005826,
  0.005753,   0.005753,    0.005753,    0.005753,
  0.005694,   0.005694,    0.005694,    0.005694,
  0.005619,   0.005619,    0.005619,    0.005619,
  0.005531,   0.005531,    0.005531,    0.005531,
  0.005465,   0.005465,    0.005465,    0.005465,
  0.005402,   0.005402,    0.005402,    0.005402,
  0.005353,   0.005353,    0.005353,    0.005353,
  0.005304,   0.005304,    0.005304,    0.005304,
  0.005236,   0.005236,    0.005236,    0.005236,
  0.005179,   0.005179,    0.005179,    0.005179,
  0.005141,   0.005141,    0.005141,    0.005141,
  0.005107,   0.005107,    0.005107,    0.005107,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005012,   0.005012,    0.005012,    0.005012,
  0.004951,   0.004951,    0.004951,    0.004951,
  0.004936,   0.004936,    0.004936,    0.004936,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005195,   0.005195,    0.005195,    0.005195,
  0.005306,   0.005306,    0.005306,    0.005306,
  0.005258,   0.005258,    0.005258,    0.005258,
  0.005083,   0.005083,    0.005083,    0.005083,
  0.004869,   0.004869,    0.004869,    0.004869,
  0.004607,   0.004607,    0.004607,    0.004607,
  0.004358,   0.004358,    0.004358,    0.004358,
  0.00401,    0.00401,     0.00401,     0.00401,
  0.003719,   0.003719,    0.003719,    0.003719,
  0.003618,   0.003618,    0.003618,    0.003618,
  0.00367,    0.00367,     0.00367,     0.00367,
  0.003765,   0.003765,    0.003765,    0.003765,
  0.003785,   0.003785,    0.003785,    0.003785,
  0.003764,   0.003764,    0.003764,    0.003764,
  0.003522,   0.003522,    0.003522,    0.003522,
  0.003267,   0.003267,    0.003267,    0.003267,
  0.003307,   0.003307,    0.003307,    0.003307,
  0.003475,   0.003475,    0.003475,    0.003475,
  0.003793,   0.003793,    0.003793,    0.003793,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004502,   0.004502,    0.004502,    0.004502,
  0.005332,   0.005332,    0.005332,    0.005332,
  0.005921,   0.005921,    0.005921,    0.005921,
  0.006096,   0.006096,    0.006096,    0.006096,
  0.006099,   0.006099,    0.006099,    0.006099,
  0.006043,   0.006043,    0.006043,    0.006043,
  0.005929,   0.005929,    0.005929,    0.005929,
  0.005722,   0.005722,    0.005722,    0.005722,
  0.005495,   0.005495,    0.005495,    0.005495,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004744,   0.004744,    0.004744,    0.004744,
  0.004714,   0.004714,    0.004714,    0.004714,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.005561,   0.005561,    0.005561,    0.005561,
  0.0056,     0.0056,      0.0056,      0.0056,
  0.005481,   0.005481,    0.005481,    0.005481,
  0.005428,   0.005428,    0.005428,    0.005428,
  0.005397,   0.005397,    0.005397,    0.005397,
  0.005323,   0.005323,    0.005323,    0.005323,
  0.005267,   0.005267,    0.005267,    0.005267,
  0.005189,   0.005189,    0.005189,    0.005189,
  0.005147,   0.005147,    0.005147,    0.005147,
  0.005173,   0.005173,    0.005173,    0.005173,
  0.005171,   0.005171,    0.005171,    0.005171,
  0.005158,   0.005158,    0.005158,    0.005158,
  0.005135,   0.005135,    0.005135,    0.005135,
  0.00508,    0.00508,     0.00508,     0.00508,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005012,   0.005012,    0.005012,    0.005012,
  0.004965,   0.004965,    0.004965,    0.004965,
  0.00492,    0.00492,     0.00492,     0.00492,
  0.004936,   0.004936,    0.004936,    0.004936,
  0.004967,   0.004967,    0.004967,    0.004967,
  0.004967,   0.004967,    0.004967,    0.004967,
  0.004967,   0.004967,    0.004967,    0.004967,
  0.004967,   0.004967,    0.004967,    0.004967,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004877,   0.004877,    0.004877,    0.004877,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004788,   0.004788,    0.004788,    0.004788,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004714,   0.004714,    0.004714,    0.004714,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004642,   0.004642,    0.004642,    0.004642,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004599,   0.004599,    0.004599,    0.004599,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.004472,   0.004472,    0.004472,    0.004472,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004628,   0.004628,    0.004628,    0.004628,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004908,   0.004908,    0.004908,    0.004908,
  0.005141,   0.005141,    0.005141,    0.005141,
  0.005307,   0.005307,    0.005307,    0.005307,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005299,   0.005299,    0.005299,    0.005299,
  0.005298,   0.005298,    0.005298,    0.005298,
  0.005339,   0.005339,    0.005339,    0.005339,
  0.005305,   0.005305,    0.005305,    0.005305,
  0.005325,   0.005325,    0.005325,    0.005325,
  0.005374,   0.005374,    0.005374,    0.005374,
  0.005416,   0.005416,    0.005416,    0.005416,
  0.005464,   0.005464,    0.005464,    0.005464,
  0.005666,   0.005666,    0.005666,    0.005666,
  0.005822,   0.005822,    0.005822,    0.005822,
  0.005839,   0.005839,    0.005839,    0.005839,
  0.00591,    0.00591,     0.00591,     0.00591,
  0.005947,   0.005947,    0.005947,    0.005947,
  0.005908,   0.005908,    0.005908,    0.005908,
  0.005895,   0.005895,    0.005895,    0.005895,
  0.005928,   0.005928,    0.005928,    0.005928,
  0.005945,   0.005945,    0.005945,    0.005945,
  0.005936,   0.005936,    0.005936,    0.005936,
  0.005843,   0.005843,    0.005843,    0.005843,
  0.005774,   0.005774,    0.005774,    0.005774,
  0.005813,   0.005813,    0.005813,    0.005813,
  0.00583,    0.00583,     0.00583,     0.00583,
  0.005767,   0.005767,    0.005767,    0.005767,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005739,   0.005739,    0.005739,    0.005739,
  0.005704,   0.005704,    0.005704,    0.005704,
  0.005626,   0.005626,    0.005626,    0.005626,
  0.005602,   0.005602,    0.005602,    0.005602,
  0.005634,   0.005634,    0.005634,    0.005634,
  0.005721,   0.005721,    0.005721,    0.005721,
  0.00583,    0.00583,     0.00583,     0.00583,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005965,   0.005965,    0.005965,    0.005965,
  0.005971,   0.005971,    0.005971,    0.005971,
  0.006008,   0.006008,    0.006008,    0.006008,
  0.006002,   0.006002,    0.006002,    0.006002,
  0.00592,    0.00592,     0.00592,     0.00592,
  0.005826,   0.005826,    0.005826,    0.005826,
  0.005822,   0.005822,    0.005822,    0.005822,
  0.005875,   0.005875,    0.005875,    0.005875,
  0.00598,    0.00598,     0.00598,     0.00598,
  0.006109,   0.006109,    0.006109,    0.006109,
  0.006149,   0.006149,    0.006149,    0.006149,
  0.006192,   0.006192,    0.006192,    0.006192,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.005963,   0.005963,    0.005963,    0.005963,
  0.005858,   0.005858,    0.005858,    0.005858,
  0.005658,   0.005658,    0.005658,    0.005658,
  0.005381,   0.005381,    0.005381,    0.005381,
  0.005333,   0.005333,    0.005333,    0.005333,
  0.005497,   0.005497,    0.005497,    0.005497,
  0.005579,   0.005579,    0.005579,    0.005579,
  0.005523,   0.005523,    0.005523,    0.005523,
  0.005624,   0.005624,    0.005624,    0.005624,
  0.005824,   0.005824,    0.005824,    0.005824,
  0.005906,   0.005906,    0.005906,    0.005906,
  0.005958,   0.005958,    0.005958,    0.005958,
  0.006056,   0.006056,    0.006056,    0.006056,
  0.006115,   0.006115,    0.006115,    0.006115,
  0.006199,   0.006199,    0.006199,    0.006199,
  0.006305,   0.006305,    0.006305,    0.006305,
  0.006307,   0.006307,    0.006307,    0.006307,
  0.006217,   0.006217,    0.006217,    0.006217,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.005661,   0.005661,    0.005661,    0.005661,
  0.005339,   0.005339,    0.005339,    0.005339,
  0.005307,   0.005307,    0.005307,    0.005307,
  0.005383,   0.005383,    0.005383,    0.005383,
  0.005458,   0.005458,    0.005458,    0.005458,
  0.00549,    0.00549,     0.00549,     0.00549,
  0.00549,    0.00549,     0.00549,     0.00549,
  0.005471,   0.005471,    0.005471,    0.005471,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005465,   0.005465,    0.005465,    0.005465,
  0.005435,   0.005435,    0.005435,    0.005435,
  0.005474,   0.005474,    0.005474,    0.005474,
  0.005519,   0.005519,    0.005519,    0.005519,
  0.005501,   0.005501,    0.005501,    0.005501,
  0.005514,   0.005514,    0.005514,    0.005514,
  0.005541,   0.005541,    0.005541,    0.005541,
  0.005573,   0.005573,    0.005573,    0.005573,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005622,   0.005622,    0.005622,    0.005622,
  0.005672,   0.005672,    0.005672,    0.005672,
  0.005708,   0.005708,    0.005708,    0.005708,
  0.005745,   0.005745,    0.005745,    0.005745,
  0.005782,   0.005782,    0.005782,    0.005782,
  0.005837,   0.005837,    0.005837,    0.005837,
  0.005912,   0.005912,    0.005912,    0.005912,
  0.005987,   0.005987,    0.005987,    0.005987,
  0.006044,   0.006044,    0.006044,    0.006044,
  0.006095,   0.006095,    0.006095,    0.006095,
  0.006183,   0.006183,    0.006183,    0.006183,
  0.006283,   0.006283,    0.006283,    0.006283,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006403,   0.006403,    0.006403,    0.006403,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.006557,   0.006557,    0.006557,    0.006557,
  0.006616,   0.006616,    0.006616,    0.006616,
  0.006636,   0.006636,    0.006636,    0.006636,
  0.006675,   0.006675,    0.006675,    0.006675,
  0.006663,   0.006663,    0.006663,    0.006663,
  0.006581,   0.006581,    0.006581,    0.006581,
  0.006549,   0.006549,    0.006549,    0.006549,
  0.006537,   0.006537,    0.006537,    0.006537,
  0.006546,   0.006546,    0.006546,    0.006546,
  0.006534,   0.006534,    0.006534,    0.006534,
  0.006503,   0.006503,    0.006503,    0.006503,
  0.006503,   0.006503,    0.006503,    0.006503,
  0.006534,   0.006534,    0.006534,    0.006534,
  0.006526,   0.006526,    0.006526,    0.006526,
  0.006471,   0.006471,    0.006471,    0.006471,
  0.006436,   0.006436,    0.006436,    0.006436,
  0.006417,   0.006417,    0.006417,    0.006417,
  0.006398,   0.006398,    0.006398,    0.006398,
  0.006378,   0.006378,    0.006378,    0.006378,
  0.006398,   0.006398,    0.006398,    0.006398,
  0.006347,   0.006347,    0.006347,    0.006347,
  0.006252,   0.006252,    0.006252,    0.006252,
  0.006208,   0.006208,    0.006208,    0.006208,
  0.006195,   0.006195,    0.006195,    0.006195,
  0.006208,   0.006208,    0.006208,    0.006208,
  0.006208,   0.006208,    0.006208,    0.006208,
  0.00622,    0.00622,     0.00622,     0.00622,
  0.006246,   0.006246,    0.006246,    0.006246,
  0.006233,   0.006233,    0.006233,    0.006233,
  0.006195,   0.006195,    0.006195,    0.006195,
  0.006176,   0.006176,    0.006176,    0.006176,
  0.006132,   0.006132,    0.006132,    0.006132,
  0.006107,   0.006107,    0.006107,    0.006107,
  0.006126,   0.006126,    0.006126,    0.006126,
  0.006107,   0.006107,    0.006107,    0.006107,
  0.006139,   0.006139,    0.006139,    0.006139,
  0.006209,   0.006209,    0.006209,    0.006209,
  0.006247,   0.006247,    0.006247,    0.006247,
  0.006231,   0.006231,    0.006231,    0.006231,
  0.00618,    0.00618,     0.00618,     0.00618,
  0.006111,   0.006111,    0.006111,    0.006111,
  0.006014,   0.006014,    0.006014,    0.006014,
  0.00597,    0.00597,     0.00597,     0.00597,
  0.006042,   0.006042,    0.006042,    0.006042,
  0.006146,   0.006146,    0.006146,    0.006146,
  0.006369,   0.006369,    0.006369,    0.006369,
  0.006578,   0.006578,    0.006578,    0.006578,
  0.006577,   0.006577,    0.006577,    0.006577,
  0.006557,   0.006557,    0.006557,    0.006557,
  0.006596,   0.006596,    0.006596,    0.006596,
  0.006675,   0.006675,    0.006675,    0.006675,
  0.006755,   0.006755,    0.006755,    0.006755,
  0.006815,   0.006815,    0.006815,    0.006815,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006896,   0.006896,    0.006896,    0.006896,
  0.006896,   0.006896,    0.006896,    0.006896,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006835,   0.006835,    0.006835,    0.006835,
  0.006815,   0.006815,    0.006815,    0.006815,
  0.006795,   0.006795,    0.006795,    0.006795,
  0.006815,   0.006815,    0.006815,    0.006815,
  0.006815,   0.006815,    0.006815,    0.006815,
  0.006795,   0.006795,    0.006795,    0.006795,
  0.006775,   0.006775,    0.006775,    0.006775,
  0.006755,   0.006755,    0.006755,    0.006755,
  0.006755,   0.006755,    0.006755,    0.006755,
  0.006755,   0.006755,    0.006755,    0.006755,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006617,   0.006617,    0.006617,    0.006617,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.006403,   0.006403,    0.006403,    0.006403,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006234,   0.006234,    0.006234,    0.006234,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.006086,   0.006086,    0.006086,    0.006086,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.006086,   0.006086,    0.006086,    0.006086,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.006215,   0.006215,    0.006215,    0.006215,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006442,   0.006442,    0.006442,    0.006442,
  0.006577,   0.006577,    0.006577,    0.006577,
  0.006775,   0.006775,    0.006775,    0.006775,
  0.006937,   0.006937,    0.006937,    0.006937,
  0.007019,   0.007019,    0.007019,    0.007019,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.007019,   0.007019,    0.007019,    0.007019,
  0.006978,   0.006978,    0.006978,    0.006978,
  0.006998,   0.006998,    0.006998,    0.006998,
  0.007039,   0.007039,    0.007039,    0.007039,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.006884,   0.006884,    0.006884,    0.006884,
  0.006531,   0.006531,    0.006531,    0.006531,
  0.006325,   0.006325,    0.006325,    0.006325,
  0.006242,   0.006242,    0.006242,    0.006242,
  0.006211,   0.006211,    0.006211,    0.006211,
  0.006191,   0.006191,    0.006191,    0.006191,
  0.006128,   0.006128,    0.006128,    0.006128,
  0.006085,   0.006085,    0.006085,    0.006085,
  0.006116,   0.006116,    0.006116,    0.006116,
  0.006148,   0.006148,    0.006148,    0.006148,
  0.006136,   0.006136,    0.006136,    0.006136,
  0.006116,   0.006116,    0.006116,    0.006116,
  0.006193,   0.006193,    0.006193,    0.006193,
  0.00634,    0.00634,     0.00634,     0.00634,
  0.006429,   0.006429,    0.006429,    0.006429,
  0.006463,   0.006463,    0.006463,    0.006463,
  0.00651,    0.00651,     0.00651,     0.00651,
  0.006555,   0.006555,    0.006555,    0.006555,
  0.006572,   0.006572,    0.006572,    0.006572,
  0.006551,   0.006551,    0.006551,    0.006551,
  0.006511,   0.006511,    0.006511,    0.006511,
  0.006494,   0.006494,    0.006494,    0.006494,
  0.006466,   0.006466,    0.006466,    0.006466,
  0.006376,   0.006376,    0.006376,    0.006376,
  0.006298,   0.006298,    0.006298,    0.006298,
  0.006253,   0.006253,    0.006253,    0.006253,
  0.006208,   0.006208,    0.006208,    0.006208,
  0.006164,   0.006164,    0.006164,    0.006164,
  0.006071,   0.006071,    0.006071,    0.006071,
  0.006028,   0.006028,    0.006028,    0.006028,
  0.005997,   0.005997,    0.005997,    0.005997,
  0.005982,   0.005982,    0.005982,    0.005982,
  0.006,      0.006,       0.006,       0.006,
  0.005919,   0.005919,    0.005919,    0.005919,
  0.005743,   0.005743,    0.005743,    0.005743,
  0.005573,   0.005573,    0.005573,    0.005573,
  0.005486,   0.005486,    0.005486,    0.005486,
  0.005435,   0.005435,    0.005435,    0.005435,
  0.005397,   0.005397,    0.005397,    0.005397,
  0.005395,   0.005395,    0.005395,    0.005395,
  0.005381,   0.005381,    0.005381,    0.005381,
  0.005296,   0.005296,    0.005296,    0.005296,
  0.005223,   0.005223,    0.005223,    0.005223,
  0.005286,   0.005286,    0.005286,    0.005286,
  0.005402,   0.005402,    0.005402,    0.005402,
  0.005391,   0.005391,    0.005391,    0.005391,
  0.005402,   0.005402,    0.005402,    0.005402,
  0.005458,   0.005458,    0.005458,    0.005458,
  0.005412,   0.005412,    0.005412,    0.005412,
  0.00538,    0.00538,     0.00538,     0.00538,
  0.00539,    0.00539,     0.00539,     0.00539,
  0.005359,   0.005359,    0.005359,    0.005359,
  0.005277,   0.005277,    0.005277,    0.005277,
  0.005196,   0.005196,    0.005196,    0.005196,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005001,   0.005001,    0.005001,    0.005001,
  0.004947,   0.004947,    0.004947,    0.004947,
  0.004895,   0.004895,    0.004895,    0.004895,
  0.004858,   0.004858,    0.004858,    0.004858,
  0.004839,   0.004839,    0.004839,    0.004839,
  0.004823,   0.004823,    0.004823,    0.004823,
  0.004793,   0.004793,    0.004793,    0.004793,
  0.004748,   0.004748,    0.004748,    0.004748,
  0.004719,   0.004719,    0.004719,    0.004719,
  0.004721,   0.004721,    0.004721,    0.004721,
  0.004691,   0.004691,    0.004691,    0.004691,
  0.004678,   0.004678,    0.004678,    0.004678,
  0.004739,   0.004739,    0.004739,    0.004739,
  0.004797,   0.004797,    0.004797,    0.004797,
  0.00478,    0.00478,     0.00478,     0.00478,
  0.004762,   0.004762,    0.004762,    0.004762,
  0.004792,   0.004792,    0.004792,    0.004792,
  0.004792,   0.004792,    0.004792,    0.004792,
  0.004807,   0.004807,    0.004807,    0.004807,
  0.00487,    0.00487,     0.00487,     0.00487,
  0.004949,   0.004949,    0.004949,    0.004949,
  0.005045,   0.005045,    0.005045,    0.005045,
  0.005111,   0.005111,    0.005111,    0.005111,
  0.005179,   0.005179,    0.005179,    0.005179,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005385,   0.005385,    0.005385,    0.005385,
  0.005598,   0.005598,    0.005598,    0.005598,
  0.00584,    0.00584,     0.00584,     0.00584,
  0.006102,   0.006102,    0.006102,    0.006102,
  0.00631,    0.00631,     0.00631,     0.00631,
  0.006435,   0.006435,    0.006435,    0.006435,
  0.006572,   0.006572,    0.006572,    0.006572,
  0.006631,   0.006631,    0.006631,    0.006631,
  0.006449,   0.006449,    0.006449,    0.006449,
  0.006233,   0.006233,    0.006233,    0.006233,
  0.006158,   0.006158,    0.006158,    0.006158,
  0.005987,   0.005987,    0.005987,    0.005987,
  0.005716,   0.005716,    0.005716,    0.005716,
  0.005666,   0.005666,    0.005666,    0.005666,
  0.005809,   0.005809,    0.005809,    0.005809,
  0.005897,   0.005897,    0.005897,    0.005897,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.005588,   0.005588,    0.005588,    0.005588,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005202,   0.005202,    0.005202,    0.005202,
  0.005284,   0.005284,    0.005284,    0.005284,
  0.005332,   0.005332,    0.005332,    0.005332,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.005479,   0.005479,    0.005479,    0.005479,
  0.005503,   0.005503,    0.005503,    0.005503,
  0.005496,   0.005496,    0.005496,    0.005496,
  0.005437,   0.005437,    0.005437,    0.005437,
  0.005431,   0.005431,    0.005431,    0.005431,
  0.005471,   0.005471,    0.005471,    0.005471,
  0.005502,   0.005502,    0.005502,    0.005502,
  0.005539,   0.005539,    0.005539,    0.005539,
  0.005554,   0.005554,    0.005554,    0.005554,
  0.005546,   0.005546,    0.005546,    0.005546,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.00551,    0.00551,     0.00551,     0.00551,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.00568,    0.00568,     0.00568,     0.00568,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005748,   0.005748,    0.005748,    0.005748,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005748,   0.005748,    0.005748,    0.005748,
  0.00584,    0.00584,     0.00584,     0.00584,
  0.005906,   0.005906,    0.005906,    0.005906,
  0.005871,   0.005871,    0.005871,    0.005871,
  0.005871,   0.005871,    0.005871,    0.005871,
  0.005839,   0.005839,    0.005839,    0.005839,
  0.005636,   0.005636,    0.005636,    0.005636,
  0.005395,   0.005395,    0.005395,    0.005395,
  0.005121,   0.005121,    0.005121,    0.005121,
  0.004844,   0.004844,    0.004844,    0.004844,
  0.004723,   0.004723,    0.004723,    0.004723,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004726,   0.004726,    0.004726,    0.004726,
  0.004526,   0.004526,    0.004526,    0.004526,
  0.00432,    0.00432,     0.00432,     0.00432,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004136,   0.004136,    0.004136,    0.004136,
  0.004028,   0.004028,    0.004028,    0.004028,
  0.003983,   0.003983,    0.003983,    0.003983,
  0.003908,   0.003908,    0.003908,    0.003908,
  0.003832,   0.003832,    0.003832,    0.003832,
  0.003789,   0.003789,    0.003789,    0.003789,
  0.003746,   0.003746,    0.003746,    0.003746,
  0.003794,   0.003794,    0.003794,    0.003794,
  0.003875,   0.003875,    0.003875,    0.003875,
  0.003846,   0.003846,    0.003846,    0.003846,
  0.003818,   0.003818,    0.003818,    0.003818,
  0.003741,   0.003741,    0.003741,    0.003741,
  0.003632,   0.003632,    0.003632,    0.003632,
  0.003636,   0.003636,    0.003636,    0.003636,
  0.003703,   0.003703,    0.003703,    0.003703,
  0.003769,   0.003769,    0.003769,    0.003769,
  0.003791,   0.003791,    0.003791,    0.003791,
  0.003764,   0.003764,    0.003764,    0.003764,
  0.003737,   0.003737,    0.003737,    0.003737,
  0.003728,   0.003728,    0.003728,    0.003728,
  0.003701,   0.003701,    0.003701,    0.003701,
  0.003675,   0.003675,    0.003675,    0.003675,
  0.003654,   0.003654,    0.003654,    0.003654,
  0.00369,    0.00369,     0.00369,     0.00369,
  0.003703,   0.003703,    0.003703,    0.003703,
  0.003659,   0.003659,    0.003659,    0.003659,
  0.003604,   0.003604,    0.003604,    0.003604,
  0.003549,   0.003549,    0.003549,    0.003549,
  0.003479,   0.003479,    0.003479,    0.003479,
  0.003468,   0.003468,    0.003468,    0.003468,
  0.003557,   0.003557,    0.003557,    0.003557,
  0.003595,   0.003595,    0.003595,    0.003595,
  0.003635,   0.003635,    0.003635,    0.003635,
  0.003661,   0.003661,    0.003661,    0.003661,
  0.003563,   0.003563,    0.003563,    0.003563,
  0.00358,    0.00358,     0.00358,     0.00358,
  0.003614,   0.003614,    0.003614,    0.003614,
  0.003676,   0.003676,    0.003676,    0.003676,
  0.003911,   0.003911,    0.003911,    0.003911,
  0.004099,   0.004099,    0.004099,    0.004099,
  0.004133,   0.004133,    0.004133,    0.004133,
  0.004136,   0.004136,    0.004136,    0.004136,
  0.004248,   0.004248,    0.004248,    0.004248,
  0.004471,   0.004471,    0.004471,    0.004471,
  0.004799,   0.004799,    0.004799,    0.004799,
  0.004999,   0.004999,    0.004999,    0.004999,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005186,   0.005186,    0.005186,    0.005186,
  0.005234,   0.005234,    0.005234,    0.005234,
  0.005218,   0.005218,    0.005218,    0.005218,
  0.005124,   0.005124,    0.005124,    0.005124,
  0.005076,   0.005076,    0.005076,    0.005076,
  0.005092,   0.005092,    0.005092,    0.005092,
  0.005092,   0.005092,    0.005092,    0.005092,
  0.005076,   0.005076,    0.005076,    0.005076,
  0.005107,   0.005107,    0.005107,    0.005107,
  0.005171,   0.005171,    0.005171,    0.005171,
  0.005154,   0.005154,    0.005154,    0.005154,
  0.005028,   0.005028,    0.005028,    0.005028,
  0.004874,   0.004874,    0.004874,    0.004874,
  0.004829,   0.004829,    0.004829,    0.004829,
  0.004874,   0.004874,    0.004874,    0.004874,
  0.00492,    0.00492,     0.00492,     0.00492,
  0.004934,   0.004934,    0.004934,    0.004934,
  0.004902,   0.004902,    0.004902,    0.004902,
  0.004871,   0.004871,    0.004871,    0.004871,
  0.004808,   0.004808,    0.004808,    0.004808,
  0.004715,   0.004715,    0.004715,    0.004715,
  0.004619,   0.004619,    0.004619,    0.004619,
  0.004556,   0.004556,    0.004556,    0.004556,
  0.00454,    0.00454,     0.00454,     0.00454,
  0.004589,   0.004589,    0.004589,    0.004589,
  0.004595,   0.004595,    0.004595,    0.004595,
  0.00458,    0.00458,     0.00458,     0.00458,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004761,   0.004761,    0.004761,    0.004761,
  0.004745,   0.004745,    0.004745,    0.004745,
  0.004716,   0.004716,    0.004716,    0.004716,
  0.004675,   0.004675,    0.004675,    0.004675,
  0.004603,   0.004603,    0.004603,    0.004603,
  0.004586,   0.004586,    0.004586,    0.004586,
  0.004632,   0.004632,    0.004632,    0.004632,
  0.00462,    0.00462,     0.00462,     0.00462,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.00444,    0.00444,     0.00444,     0.00444,
  0.004387,   0.004387,    0.004387,    0.004387,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004412,   0.004412,    0.004412,    0.004412,
  0.004402,   0.004402,    0.004402,    0.004402,
  0.004016,   0.004016,    0.004016,    0.004016,
  0.003905,   0.003905,    0.003905,    0.003905,
  0.004067,   0.004067,    0.004067,    0.004067,
  0.004219,   0.004219,    0.004219,    0.004219,
  0.004369,   0.004369,    0.004369,    0.004369,
  0.004479,   0.004479,    0.004479,    0.004479,
  0.004465,   0.004465,    0.004465,    0.004465,
  0.004383,   0.004383,    0.004383,    0.004383,
  0.00424,    0.00424,     0.00424,     0.00424,
  0.004118,   0.004118,    0.004118,    0.004118,
  0.004083,   0.004083,    0.004083,    0.004083,
  0.004032,   0.004032,    0.004032,    0.004032,
  0.003942,   0.003942,    0.003942,    0.003942,
  0.003846,   0.003846,    0.003846,    0.003846,
  0.003722,   0.003722,    0.003722,    0.003722,
  0.003651,   0.003651,    0.003651,    0.003651,
  0.003644,   0.003644,    0.003644,    0.003644,
  0.003625,   0.003625,    0.003625,    0.003625,
  0.003644,   0.003644,    0.003644,    0.003644,
  0.003657,   0.003657,    0.003657,    0.003657,
  0.00358,    0.00358,     0.00358,     0.00358,
  0.003582,   0.003582,    0.003582,    0.003582,
  0.003681,   0.003681,    0.003681,    0.003681,
  0.003677,   0.003677,    0.003677,    0.003677,
  0.00363,    0.00363,     0.00363,     0.00363,
  0.003615,   0.003615,    0.003615,    0.003615,
  0.0036,     0.0036,      0.0036,      0.0036,
  0.003543,   0.003543,    0.003543,    0.003543,
  0.003443,   0.003443,    0.003443,    0.003443,
  0.003443,   0.003443,    0.003443,    0.003443,
  0.00352,    0.00352,     0.00352,     0.00352,
  0.003412,   0.003412,    0.003412,    0.003412,
  0.003281,   0.003281,    0.003281,    0.003281,
  0.003345,   0.003345,    0.003345,    0.003345,
  0.003488,   0.003488,    0.003488,    0.003488,
  0.003639,   0.003639,    0.003639,    0.003639,
  0.003868,   0.003868,    0.003868,    0.003868,
  0.004059,   0.004059,    0.004059,    0.004059,
  0.004073,   0.004073,    0.004073,    0.004073,
  0.003973,   0.003973,    0.003973,    0.003973,
  0.003847,   0.003847,    0.003847,    0.003847,
  0.003755,   0.003755,    0.003755,    0.003755,
  0.003728,   0.003728,    0.003728,    0.003728,
  0.003702,   0.003702,    0.003702,    0.003702,
  0.003501,   0.003501,    0.003501,    0.003501,
  0.003324,   0.003324,    0.003324,    0.003324,
  0.003302,   0.003302,    0.003302,    0.003302,
  0.003247,   0.003247,    0.003247,    0.003247,
  0.003183,   0.003183,    0.003183,    0.003183,
  0.003175,   0.003175,    0.003175,    0.003175,
  0.00318,    0.00318,     0.00318,     0.00318,
  0.003186,   0.003186,    0.003186,    0.003186,
  0.003217,   0.003217,    0.003217,    0.003217,
  0.003188,   0.003188,    0.003188,    0.003188,
  0.003139,   0.003139,    0.003139,    0.003139,
  0.003149,   0.003149,    0.003149,    0.003149,
  0.003198,   0.003198,    0.003198,    0.003198,
  0.003333,   0.003333,    0.003333,    0.003333,
  0.003501,   0.003501,    0.003501,    0.003501,
  0.003564,   0.003564,    0.003564,    0.003564,
  0.003595,   0.003595,    0.003595,    0.003595,
  0.003626,   0.003626,    0.003626,    0.003626,
  0.003626,   0.003626,    0.003626,    0.003626,
  0.003673,   0.003673,    0.003673,    0.003673,
  0.003689,   0.003689,    0.003689,    0.003689,
  0.003657,   0.003657,    0.003657,    0.003657,
  0.003657,   0.003657,    0.003657,    0.003657,
  0.003673,   0.003673,    0.003673,    0.003673,
  0.003642,   0.003642,    0.003642,    0.003642,
  0.003595,   0.003595,    0.003595,    0.003595,
  0.003579,   0.003579,    0.003579,    0.003579,
  0.003626,   0.003626,    0.003626,    0.003626,
  0.00369,    0.00369,     0.00369,     0.00369,
  0.003658,   0.003658,    0.003658,    0.003658,
  0.003595,   0.003595,    0.003595,    0.003595,
  0.003627,   0.003627,    0.003627,    0.003627,
  0.003674,   0.003674,    0.003674,    0.003674,
  0.003736,   0.003736,    0.003736,    0.003736,
  0.003846,   0.003846,    0.003846,    0.003846,
  0.003925,   0.003925,    0.003925,    0.003925,
  0.004067,   0.004067,    0.004067,    0.004067,
  0.004352,   0.004352,    0.004352,    0.004352,
  0.004526,   0.004526,    0.004526,    0.004526,
  0.00454,    0.00454,     0.00454,     0.00454,
  0.004429,   0.004429,    0.004429,    0.004429,
  0.004256,   0.004256,    0.004256,    0.004256,
  0.004303,   0.004303,    0.004303,    0.004303,
  0.004461,   0.004461,    0.004461,    0.004461,
  0.004555,   0.004555,    0.004555,    0.004555,
  0.004634,   0.004634,    0.004634,    0.004634,
  0.004761,   0.004761,    0.004761,    0.004761,
  0.004887,   0.004887,    0.004887,    0.004887,
  0.004965,   0.004965,    0.004965,    0.004965,
  0.005012,   0.005012,    0.005012,    0.005012,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.00517,    0.00517,     0.00517,     0.00517,
  0.005187,   0.005187,    0.005187,    0.005187,
  0.005203,   0.005203,    0.005203,    0.005203,
  0.005267,   0.005267,    0.005267,    0.005267,
  0.005363,   0.005363,    0.005363,    0.005363,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.00551,    0.00551,     0.00551,     0.00551,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.005444,   0.005444,    0.005444,    0.005444,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005498,   0.005498,    0.005498,    0.005498,
  0.005456,   0.005456,    0.005456,    0.005456,
  0.005448,   0.005448,    0.005448,    0.005448,
  0.005423,   0.005423,    0.005423,    0.005423,
  0.00543,    0.00543,     0.00543,     0.00543,
  0.005424,   0.005424,    0.005424,    0.005424,
  0.005402,   0.005402,    0.005402,    0.005402,
  0.005407,   0.005407,    0.005407,    0.005407,
  0.005407,   0.005407,    0.005407,    0.005407,
  0.00547,    0.00547,     0.00547,     0.00547,
  0.005519,   0.005519,    0.005519,    0.005519,
  0.005519,   0.005519,    0.005519,    0.005519,
  0.005465,   0.005465,    0.005465,    0.005465,
  0.005424,   0.005424,    0.005424,    0.005424,
  0.005465,   0.005465,    0.005465,    0.005465,
  0.005448,   0.005448,    0.005448,    0.005448,
  0.005367,   0.005367,    0.005367,    0.005367,
  0.00544,    0.00544,     0.00544,     0.00544,
  0.0055,     0.0055,      0.0055,      0.0055,
  0.005494,   0.005494,    0.005494,    0.005494,
  0.005551,   0.005551,    0.005551,    0.005551,
  0.005597,   0.005597,    0.005597,    0.005597,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.00551,    0.00551,     0.00551,     0.00551,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.00551,    0.00551,     0.00551,     0.00551,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005444,   0.005444,    0.005444,    0.005444,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005697,   0.005697,    0.005697,    0.005697,
  0.005755,   0.005755,    0.005755,    0.005755,
  0.005767,   0.005767,    0.005767,    0.005767,
  0.00578,    0.00578,     0.00578,     0.00578,
  0.005764,   0.005764,    0.005764,    0.005764,
  0.005724,   0.005724,    0.005724,    0.005724,
  0.00563,    0.00563,     0.00563,     0.00563,
  0.005484,   0.005484,    0.005484,    0.005484,
  0.005408,   0.005408,    0.005408,    0.005408,
  0.005377,   0.005377,    0.005377,    0.005377,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.00527,    0.00527,     0.00527,     0.00527,
  0.005234,   0.005234,    0.005234,    0.005234,
  0.005171,   0.005171,    0.005171,    0.005171,
  0.005195,   0.005195,    0.005195,    0.005195,
  0.005364,   0.005364,    0.005364,    0.005364,
  0.00549,    0.00549,     0.00549,     0.00549,
  0.005494,   0.005494,    0.005494,    0.005494,
  0.005511,   0.005511,    0.005511,    0.005511,
  0.005534,   0.005534,    0.005534,    0.005534,
  0.005483,   0.005483,    0.005483,    0.005483,
  0.005415,   0.005415,    0.005415,    0.005415,
  0.005422,   0.005422,    0.005422,    0.005422,
  0.005437,   0.005437,    0.005437,    0.005437,
  0.005425,   0.005425,    0.005425,    0.005425,
  0.005405,   0.005405,    0.005405,    0.005405,
  0.00537,    0.00537,     0.00537,     0.00537,
  0.005333,   0.005333,    0.005333,    0.005333,
  0.005314,   0.005314,    0.005314,    0.005314,
  0.005249,   0.005249,    0.005249,    0.005249,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005014,   0.005014,    0.005014,    0.005014,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005249,   0.005249,    0.005249,    0.005249,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.005479,   0.005479,    0.005479,    0.005479,
  0.005495,   0.005495,    0.005495,    0.005495,
  0.005425,   0.005425,    0.005425,    0.005425,
  0.005386,   0.005386,    0.005386,    0.005386,
  0.005389,   0.005389,    0.005389,    0.005389,
  0.005471,   0.005471,    0.005471,    0.005471,
  0.005605,   0.005605,    0.005605,    0.005605,
  0.005708,   0.005708,    0.005708,    0.005708,
  0.005795,   0.005795,    0.005795,    0.005795,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.006118,   0.006118,    0.006118,    0.006118,
  0.006127,   0.006127,    0.006127,    0.006127,
  0.006077,   0.006077,    0.006077,    0.006077,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.005935,   0.005935,    0.005935,    0.005935,
  0.0059,     0.0059,      0.0059,      0.0059,
  0.005897,   0.005897,    0.005897,    0.005897,
  0.00584,    0.00584,     0.00584,     0.00584,
  0.005784,   0.005784,    0.005784,    0.005784,
  0.005736,   0.005736,    0.005736,    0.005736,
  0.005759,   0.005759,    0.005759,    0.005759,
  0.005814,   0.005814,    0.005814,    0.005814,
  0.005712,   0.005712,    0.005712,    0.005712,
  0.005617,   0.005617,    0.005617,    0.005617,
  0.005681,   0.005681,    0.005681,    0.005681,
  0.006097,   0.006097,    0.006097,    0.006097,
  0.006654,   0.006654,    0.006654,    0.006654,
  0.006924,   0.006924,    0.006924,    0.006924,
  0.006998,   0.006998,    0.006998,    0.006998,
  0.00704,    0.00704,     0.00704,     0.00704,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007186,   0.007186,    0.007186,    0.007186,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007239,   0.007239,    0.007239,    0.007239,
  0.007272,   0.007272,    0.007272,    0.007272,
  0.007284,   0.007284,    0.007284,    0.007284,
  0.007156,   0.007156,    0.007156,    0.007156,
  0.006976,   0.006976,    0.006976,    0.006976,
  0.00683,    0.00683,     0.00683,     0.00683,
  0.006718,   0.006718,    0.006718,    0.006718,
  0.006558,   0.006558,    0.006558,    0.006558,
  0.006352,   0.006352,    0.006352,    0.006352,
  0.005805,   0.005805,    0.005805,    0.005805,
  0.005242,   0.005242,    0.005242,    0.005242,
  0.005031,   0.005031,    0.005031,    0.005031,
  0.004872,   0.004872,    0.004872,    0.004872,
  0.004785,   0.004785,    0.004785,    0.004785,
  0.004777,   0.004777,    0.004777,    0.004777,
  0.004889,   0.004889,    0.004889,    0.004889,
  0.005159,   0.005159,    0.005159,    0.005159,
  0.005254,   0.005254,    0.005254,    0.005254,
  0.005057,   0.005057,    0.005057,    0.005057,
  0.004733,   0.004733,    0.004733,    0.004733,
  0.004405,   0.004405,    0.004405,    0.004405,
  0.004309,   0.004309,    0.004309,    0.004309,
  0.004307,   0.004307,    0.004307,    0.004307,
  0.004114,   0.004114,    0.004114,    0.004114,
  0.003872,   0.003872,    0.003872,    0.003872,
  0.003738,   0.003738,    0.003738,    0.003738,
  0.003579,   0.003579,    0.003579,    0.003579,
  0.003586,   0.003586,    0.003586,    0.003586,
  0.003555,   0.003555,    0.003555,    0.003555,
  0.003354,   0.003354,    0.003354,    0.003354,
  0.003389,   0.003389,    0.003389,    0.003389,
  0.003218,   0.003218,    0.003218,    0.003218,
  0.002871,   0.002871,    0.002871,    0.002871,
  0.002822,   0.002822,    0.002822,    0.002822,
  0.002759,   0.002759,    0.002759,    0.002759,
  0.002874,   0.002874,    0.002874,    0.002874,
  0.003509,   0.003509,    0.003509,    0.003509,
  0.00424,    0.00424,     0.00424,     0.00424,
  0.004759,   0.004759,    0.004759,    0.004759,
  0.00494,    0.00494,     0.00494,     0.00494,
  0.00494,    0.00494,     0.00494,     0.00494,
  0.004737,   0.004737,    0.004737,    0.004737,
  0.004767,   0.004767,    0.004767,    0.004767,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005931,   0.005931,    0.005931,    0.005931,
  0.006174,   0.006174,    0.006174,    0.006174,
  0.0063,     0.0063,      0.0063,      0.0063,
  0.006457,   0.006457,    0.006457,    0.006457,
  0.006536,   0.006536,    0.006536,    0.006536,
  0.00653,    0.00653,     0.00653,     0.00653,
  0.00653,    0.00653,     0.00653,     0.00653,
  0.00653,    0.00653,     0.00653,     0.00653,
  0.006632,   0.006632,    0.006632,    0.006632,
  0.006408,   0.006408,    0.006408,    0.006408,
  0.005689,   0.005689,    0.005689,    0.005689,
  0.005171,   0.005171,    0.005171,    0.005171,
  0.004992,   0.004992,    0.004992,    0.004992,
  0.004859,   0.004859,    0.004859,    0.004859,
  0.004723,   0.004723,    0.004723,    0.004723,
  0.004673,   0.004673,    0.004673,    0.004673,
  0.004703,   0.004703,    0.004703,    0.004703,
  0.004721,   0.004721,    0.004721,    0.004721,
  0.004744,   0.004744,    0.004744,    0.004744,
  0.004735,   0.004735,    0.004735,    0.004735,
  0.004677,   0.004677,    0.004677,    0.004677,
  0.004635,   0.004635,    0.004635,    0.004635,
  0.004621,   0.004621,    0.004621,    0.004621,
  0.004593,   0.004593,    0.004593,    0.004593,
  0.004507,   0.004507,    0.004507,    0.004507,
  0.004344,   0.004344,    0.004344,    0.004344,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004188,   0.004188,    0.004188,    0.004188,
  0.004149,   0.004149,    0.004149,    0.004149,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.00401,    0.00401,     0.00401,     0.00401,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003871,   0.003871,    0.003871,    0.003871,
  0.003936,   0.003936,    0.003936,    0.003936,
  0.003981,   0.003981,    0.003981,    0.003981,
  0.004026,   0.004026,    0.004026,    0.004026,
  0.004089,   0.004089,    0.004089,    0.004089,
  0.004049,   0.004049,    0.004049,    0.004049,
  0.003931,   0.003931,    0.003931,    0.003931,
  0.003867,   0.003867,    0.003867,    0.003867,
  0.003845,   0.003845,    0.003845,    0.003845,
  0.003827,   0.003827,    0.003827,    0.003827,
  0.003841,   0.003841,    0.003841,    0.003841,
  0.003949,   0.003949,    0.003949,    0.003949,
  0.004026,   0.004026,    0.004026,    0.004026,
  0.00404,    0.00404,     0.00404,     0.00404,
  0.004023,   0.004023,    0.004023,    0.004023,
  0.003974,   0.003974,    0.003974,    0.003974,
  0.003999,   0.003999,    0.003999,    0.003999,
  0.004005,   0.004005,    0.004005,    0.004005,
  0.004032,   0.004032,    0.004032,    0.004032,
  0.004095,   0.004095,    0.004095,    0.004095,
  0.004108,   0.004108,    0.004108,    0.004108,
  0.004152,   0.004152,    0.004152,    0.004152,
  0.004181,   0.004181,    0.004181,    0.004181,
  0.004147,   0.004147,    0.004147,    0.004147,
  0.004147,   0.004147,    0.004147,    0.004147,
  0.004225,   0.004225,    0.004225,    0.004225,
  0.004256,   0.004256,    0.004256,    0.004256,
  0.00424,    0.00424,     0.00424,     0.00424,
  0.00424,    0.00424,     0.00424,     0.00424,
  0.004288,   0.004288,    0.004288,    0.004288,
  0.004367,   0.004367,    0.004367,    0.004367,
  0.004446,   0.004446,    0.004446,    0.004446,
  0.00451,    0.00451,     0.00451,     0.00451,
  0.004574,   0.004574,    0.004574,    0.004574,
  0.004497,   0.004497,    0.004497,    0.004497,
  0.004421,   0.004421,    0.004421,    0.004421,
  0.004534,   0.004534,    0.004534,    0.004534,
  0.004569,   0.004569,    0.004569,    0.004569,
  0.004574,   0.004574,    0.004574,    0.004574,
  0.004654,   0.004654,    0.004654,    0.004654,
  0.004619,   0.004619,    0.004619,    0.004619,
  0.004426,   0.004426,    0.004426,    0.004426,
  0.004118,   0.004118,    0.004118,    0.004118,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.004211,   0.004211,    0.004211,    0.004211,
  0.004527,   0.004527,    0.004527,    0.004527,
  0.00475,    0.00475,     0.00475,     0.00475,
  0.004719,   0.004719,    0.004719,    0.004719,
  0.004584,   0.004584,    0.004584,    0.004584,
  0.004475,   0.004475,    0.004475,    0.004475,
  0.004545,   0.004545,    0.004545,    0.004545,
  0.004526,   0.004526,    0.004526,    0.004526,
  0.004425,   0.004425,    0.004425,    0.004425,
  0.0044,     0.0044,      0.0044,      0.0044,
  0.0044,     0.0044,      0.0044,      0.0044,
  0.004419,   0.004419,    0.004419,    0.004419,
  0.004533,   0.004533,    0.004533,    0.004533,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004705,   0.004705,    0.004705,    0.004705,
  0.004736,   0.004736,    0.004736,    0.004736,
  0.004835,   0.004835,    0.004835,    0.004835,
  0.004859,   0.004859,    0.004859,    0.004859,
  0.00495,    0.00495,     0.00495,     0.00495,
  0.005111,   0.005111,    0.005111,    0.005111,
  0.00508,    0.00508,     0.00508,     0.00508,
  0.004999,   0.004999,    0.004999,    0.004999,
  0.005031,   0.005031,    0.005031,    0.005031,
  0.00508,    0.00508,     0.00508,     0.00508,
  0.005136,   0.005136,    0.005136,    0.005136,
  0.005224,   0.005224,    0.005224,    0.005224,
  0.005307,   0.005307,    0.005307,    0.005307,
  0.005374,   0.005374,    0.005374,    0.005374,
  0.005368,   0.005368,    0.005368,    0.005368,
  0.005294,   0.005294,    0.005294,    0.005294,
  0.005207,   0.005207,    0.005207,    0.005207,
  0.005156,   0.005156,    0.005156,    0.005156,
  0.005139,   0.005139,    0.005139,    0.005139,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.005059,   0.005059,    0.005059,    0.005059,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005237,   0.005237,    0.005237,    0.005237,
  0.005314,   0.005314,    0.005314,    0.005314,
  0.005296,   0.005296,    0.005296,    0.005296,
  0.005114,   0.005114,    0.005114,    0.005114,
  0.004818,   0.004818,    0.004818,    0.004818,
  0.004671,   0.004671,    0.004671,    0.004671,
  0.004668,   0.004668,    0.004668,    0.004668,
  0.004593,   0.004593,    0.004593,    0.004593,
  0.004392,   0.004392,    0.004392,    0.004392,
  0.004266,   0.004266,    0.004266,    0.004266,
  0.004213,   0.004213,    0.004213,    0.004213,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.004147,   0.004147,    0.004147,    0.004147,
  0.004068,   0.004068,    0.004068,    0.004068,
  0.004106,   0.004106,    0.004106,    0.004106,
  0.004279,   0.004279,    0.004279,    0.004279,
  0.004397,   0.004397,    0.004397,    0.004397,
  0.004357,   0.004357,    0.004357,    0.004357,
  0.004311,   0.004311,    0.004311,    0.004311,
  0.004368,   0.004368,    0.004368,    0.004368,
  0.004478,   0.004478,    0.004478,    0.004478,
  0.004559,   0.004559,    0.004559,    0.004559,
  0.004584,   0.004584,    0.004584,    0.004584,
  0.004592,   0.004592,    0.004592,    0.004592,
  0.004629,   0.004629,    0.004629,    0.004629,
  0.004752,   0.004752,    0.004752,    0.004752,
  0.004863,   0.004863,    0.004863,    0.004863,
  0.004893,   0.004893,    0.004893,    0.004893,
  0.004897,   0.004897,    0.004897,    0.004897,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004919,   0.004919,    0.004919,    0.004919,
  0.004933,   0.004933,    0.004933,    0.004933,
  0.004917,   0.004917,    0.004917,    0.004917,
  0.004856,   0.004856,    0.004856,    0.004856,
  0.004768,   0.004768,    0.004768,    0.004768,
  0.004666,   0.004666,    0.004666,    0.004666,
  0.004625,   0.004625,    0.004625,    0.004625,
  0.004585,   0.004585,    0.004585,    0.004585,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.004364,   0.004364,    0.004364,    0.004364,
  0.004088,   0.004088,    0.004088,    0.004088,
  0.003873,   0.003873,    0.003873,    0.003873,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.003947,   0.003947,    0.003947,    0.003947,
  0.003824,   0.003824,    0.003824,    0.003824,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.003947,   0.003947,    0.003947,    0.003947,
  0.004152,   0.004152,    0.004152,    0.004152,
  0.00452,    0.00452,     0.00452,     0.00452,
  0.005084,   0.005084,    0.005084,    0.005084,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005003,   0.005003,    0.005003,    0.005003,
  0.004777,   0.004777,    0.004777,    0.004777,
  0.004635,   0.004635,    0.004635,    0.004635,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004473,   0.004473,    0.004473,    0.004473,
  0.004434,   0.004434,    0.004434,    0.004434,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004369,   0.004369,    0.004369,    0.004369,
  0.004327,   0.004327,    0.004327,    0.004327,
  0.004357,   0.004357,    0.004357,    0.004357,
  0.004368,   0.004368,    0.004368,    0.004368,
  0.004287,   0.004287,    0.004287,    0.004287,
  0.00418,    0.00418,     0.00418,     0.00418,
  0.004161,   0.004161,    0.004161,    0.004161,
  0.004155,   0.004155,    0.004155,    0.004155,
  0.004194,   0.004194,    0.004194,    0.004194,
  0.004258,   0.004258,    0.004258,    0.004258,
  0.004368,   0.004368,    0.004368,    0.004368,
  0.004504,   0.004504,    0.004504,    0.004504,
  0.004573,   0.004573,    0.004573,    0.004573,
  0.004616,   0.004616,    0.004616,    0.004616,
  0.004621,   0.004621,    0.004621,    0.004621,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.00457,    0.00457,     0.00457,     0.00457,
  0.004546,   0.004546,    0.004546,    0.004546,
  0.00453,    0.00453,     0.00453,     0.00453,
  0.004488,   0.004488,    0.004488,    0.004488,
  0.004455,   0.004455,    0.004455,    0.004455,
  0.004414,   0.004414,    0.004414,    0.004414,
  0.004389,   0.004389,    0.004389,    0.004389,
  0.004373,   0.004373,    0.004373,    0.004373,
  0.004336,   0.004336,    0.004336,    0.004336,
  0.004303,   0.004303,    0.004303,    0.004303,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004367,   0.004367,    0.004367,    0.004367,
  0.004383,   0.004383,    0.004383,    0.004383,
  0.00443,    0.00443,     0.00443,     0.00443,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004461,   0.004461,    0.004461,    0.004461,
  0.004493,   0.004493,    0.004493,    0.004493,
  0.004479,   0.004479,    0.004479,    0.004479,
  0.004509,   0.004509,    0.004509,    0.004509,
  0.004508,   0.004508,    0.004508,    0.004508,
  0.004524,   0.004524,    0.004524,    0.004524,
  0.004646,   0.004646,    0.004646,    0.004646,
  0.004767,   0.004767,    0.004767,    0.004767,
  0.0048,     0.0048,      0.0048,      0.0048,
  0.004578,   0.004578,    0.004578,    0.004578,
  0.004281,   0.004281,    0.004281,    0.004281,
  0.004154,   0.004154,    0.004154,    0.004154,
  0.004181,   0.004181,    0.004181,    0.004181,
  0.0042,     0.0042,      0.0042,      0.0042,
  0.004117,   0.004117,    0.004117,    0.004117,
  0.004103,   0.004103,    0.004103,    0.004103,
  0.00411,    0.00411,     0.00411,     0.00411,
  0.003978,   0.003978,    0.003978,    0.003978,
  0.003857,   0.003857,    0.003857,    0.003857,
  0.003772,   0.003772,    0.003772,    0.003772,
  0.003772,   0.003772,    0.003772,    0.003772,
  0.003866,   0.003866,    0.003866,    0.003866,
  0.00374,    0.00374,     0.00374,     0.00374,
  0.003624,   0.003624,    0.003624,    0.003624,
  0.00362,    0.00362,     0.00362,     0.00362,
  0.00357,    0.00357,     0.00357,     0.00357,
  0.003758,   0.003758,    0.003758,    0.003758,
  0.004075,   0.004075,    0.004075,    0.004075,
  0.004331,   0.004331,    0.004331,    0.004331,
  0.004579,   0.004579,    0.004579,    0.004579,
  0.004732,   0.004732,    0.004732,    0.004732,
  0.00479,    0.00479,     0.00479,     0.00479,
  0.004831,   0.004831,    0.004831,    0.004831,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004754,   0.004754,    0.004754,    0.004754,
  0.004731,   0.004731,    0.004731,    0.004731,
  0.004724,   0.004724,    0.004724,    0.004724,
  0.004704,   0.004704,    0.004704,    0.004704,
  0.00466,    0.00466,     0.00466,     0.00466,
  0.004639,   0.004639,    0.004639,    0.004639,
  0.004717,   0.004717,    0.004717,    0.004717,
  0.004748,   0.004748,    0.004748,    0.004748,
  0.004698,   0.004698,    0.004698,    0.004698,
  0.004744,   0.004744,    0.004744,    0.004744,
  0.004761,   0.004761,    0.004761,    0.004761,
  0.004672,   0.004672,    0.004672,    0.004672,
  0.004599,   0.004599,    0.004599,    0.004599,
  0.004531,   0.004531,    0.004531,    0.004531,
  0.004424,   0.004424,    0.004424,    0.004424,
  0.004291,   0.004291,    0.004291,    0.004291,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004527,   0.004527,    0.004527,    0.004527,
  0.004816,   0.004816,    0.004816,    0.004816,
  0.005096,   0.005096,    0.005096,    0.005096,
  0.005199,   0.005199,    0.005199,    0.005199,
  0.005161,   0.005161,    0.005161,    0.005161,
  0.005072,   0.005072,    0.005072,    0.005072,
  0.005066,   0.005066,    0.005066,    0.005066,
  0.005026,   0.005026,    0.005026,    0.005026,
  0.004768,   0.004768,    0.004768,    0.004768,
  0.004609,   0.004609,    0.004609,    0.004609,
  0.004631,   0.004631,    0.004631,    0.004631,
  0.004674,   0.004674,    0.004674,    0.004674,
  0.004665,   0.004665,    0.004665,    0.004665,
  0.00443,    0.00443,     0.00443,     0.00443,
  0.004076,   0.004076,    0.004076,    0.004076,
  0.003911,   0.003911,    0.003911,    0.003911,
  0.003911,   0.003911,    0.003911,    0.003911,
  0.003918,   0.003918,    0.003918,    0.003918,
  0.003926,   0.003926,    0.003926,    0.003926,
  0.003965,   0.003965,    0.003965,    0.003965,
  0.004043,   0.004043,    0.004043,    0.004043,
  0.004196,   0.004196,    0.004196,    0.004196,
  0.004392,   0.004392,    0.004392,    0.004392,
  0.004536,   0.004536,    0.004536,    0.004536,
  0.004671,   0.004671,    0.004671,    0.004671,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004972,   0.004972,    0.004972,    0.004972,
  0.005047,   0.005047,    0.005047,    0.005047,
  0.005074,   0.005074,    0.005074,    0.005074,
  0.004991,   0.004991,    0.004991,    0.004991,
  0.004875,   0.004875,    0.004875,    0.004875,
  0.004807,   0.004807,    0.004807,    0.004807,
  0.004776,   0.004776,    0.004776,    0.004776,
  0.004779,   0.004779,    0.004779,    0.004779,
  0.004796,   0.004796,    0.004796,    0.004796,
  0.004871,   0.004871,    0.004871,    0.004871,
  0.004943,   0.004943,    0.004943,    0.004943,
  0.004984,   0.004984,    0.004984,    0.004984,
  0.005,      0.005,       0.005,       0.005,
  0.005017,   0.005017,    0.005017,    0.005017,
  0.005061,   0.005061,    0.005061,    0.005061,
  0.005056,   0.005056,    0.005056,    0.005056,
  0.005012,   0.005012,    0.005012,    0.005012,
  0.004973,   0.004973,    0.004973,    0.004973,
  0.004898,   0.004898,    0.004898,    0.004898,
  0.004848,   0.004848,    0.004848,    0.004848,
  0.004886,   0.004886,    0.004886,    0.004886,
  0.004949,   0.004949,    0.004949,    0.004949,
  0.005024,   0.005024,    0.005024,    0.005024,
  0.005118,   0.005118,    0.005118,    0.005118,
  0.005272,   0.005272,    0.005272,    0.005272,
  0.005483,   0.005483,    0.005483,    0.005483,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005558,   0.005558,    0.005558,    0.005558,
  0.005369,   0.005369,    0.005369,    0.005369,
  0.005066,   0.005066,    0.005066,    0.005066,
  0.004877,   0.004877,    0.004877,    0.004877,
  0.004919,   0.004919,    0.004919,    0.004919,
  0.005017,   0.005017,    0.005017,    0.005017,
  0.005065,   0.005065,    0.005065,    0.005065,
  0.005148,   0.005148,    0.005148,    0.005148,
  0.00491,    0.00491,     0.00491,     0.00491,
  0.004351,   0.004351,    0.004351,    0.004351,
  0.003922,   0.003922,    0.003922,    0.003922,
  0.003766,   0.003766,    0.003766,    0.003766,
  0.003591,   0.003591,    0.003591,    0.003591,
  0.003305,   0.003305,    0.003305,    0.003305,
  0.003269,   0.003269,    0.003269,    0.003269,
  0.003444,   0.003444,    0.003444,    0.003444,
  0.00372,    0.00372,     0.00372,     0.00372,
  0.004249,   0.004249,    0.004249,    0.004249,
  0.004555,   0.004555,    0.004555,    0.004555,
  0.00444,    0.00444,     0.00444,     0.00444,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004116,   0.004116,    0.004116,    0.004116,
  0.004177,   0.004177,    0.004177,    0.004177,
  0.004161,   0.004161,    0.004161,    0.004161,
  0.004148,   0.004148,    0.004148,    0.004148,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004278,   0.004278,    0.004278,    0.004278,
  0.004341,   0.004341,    0.004341,    0.004341,
  0.004432,   0.004432,    0.004432,    0.004432,
  0.004383,   0.004383,    0.004383,    0.004383,
  0.004241,   0.004241,    0.004241,    0.004241,
  0.00413,    0.00413,     0.00413,     0.00413,
  0.00402,    0.00402,     0.00402,     0.00402,
  0.003926,   0.003926,    0.003926,    0.003926,
  0.003848,   0.003848,    0.003848,    0.003848,
  0.003805,   0.003805,    0.003805,    0.003805,
  0.003683,   0.003683,    0.003683,    0.003683,
  0.003383,   0.003383,    0.003383,    0.003383,
  0.003272,   0.003272,    0.003272,    0.003272,
  0.00335,    0.00335,     0.00335,     0.00335,
  0.003316,   0.003316,    0.003316,    0.003316,
  0.003313,   0.003313,    0.003313,    0.003313,
  0.003628,   0.003628,    0.003628,    0.003628,
  0.004007,   0.004007,    0.004007,    0.004007,
  0.004056,   0.004056,    0.004056,    0.004056,
  0.003858,   0.003858,    0.003858,    0.003858,
  0.003903,   0.003903,    0.003903,    0.003903,
  0.00432,    0.00432,     0.00432,     0.00432,
  0.004256,   0.004256,    0.004256,    0.004256,
  0.00383,    0.00383,     0.00383,     0.00383,
  0.003464,   0.003464,    0.003464,    0.003464,
  0.003548,   0.003548,    0.003548,    0.003548,
  0.003607,   0.003607,    0.003607,    0.003607,
  0.003247,   0.003247,    0.003247,    0.003247,
  0.003125,   0.003125,    0.003125,    0.003125,
  0.003003,   0.003003,    0.003003,    0.003003,
  0.00317,    0.00317,     0.00317,     0.00317,
  0.003344,   0.003344,    0.003344,    0.003344,
  0.003346,   0.003346,    0.003346,    0.003346,
  0.003312,   0.003312,    0.003312,    0.003312,
  0.003188,   0.003188,    0.003188,    0.003188,
  0.003262,   0.003262,    0.003262,    0.003262,
  0.003274,   0.003274,    0.003274,    0.003274,
  0.003286,   0.003286,    0.003286,    0.003286,
  0.003406,   0.003406,    0.003406,    0.003406,
  0.003484,   0.003484,    0.003484,    0.003484,
  0.003548,   0.003548,    0.003548,    0.003548,
  0.003597,   0.003597,    0.003597,    0.003597,
  0.003707,   0.003707,    0.003707,    0.003707,
  0.003835,   0.003835,    0.003835,    0.003835,
  0.003889,   0.003889,    0.003889,    0.003889,
  0.003947,   0.003947,    0.003947,    0.003947,
  0.003969,   0.003969,    0.003969,    0.003969,
  0.003826,   0.003826,    0.003826,    0.003826,
  0.003692,   0.003692,    0.003692,    0.003692,
  0.003683,   0.003683,    0.003683,    0.003683,
  0.003678,   0.003678,    0.003678,    0.003678,
  0.003708,   0.003708,    0.003708,    0.003708,
  0.003722,   0.003722,    0.003722,    0.003722,
  0.003658,   0.003658,    0.003658,    0.003658,
  0.003626,   0.003626,    0.003626,    0.003626,
  0.003673,   0.003673,    0.003673,    0.003673,
  0.003972,   0.003972,    0.003972,    0.003972,
  0.004476,   0.004476,    0.004476,    0.004476,
  0.004886,   0.004886,    0.004886,    0.004886,
  0.005235,   0.005235,    0.005235,    0.005235,
  0.005545,   0.005545,    0.005545,    0.005545,
  0.00582,    0.00582,     0.00582,     0.00582,
  0.006106,   0.006106,    0.006106,    0.006106,
  0.00629,    0.00629,     0.00629,     0.00629,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006403,   0.006403,    0.006403,    0.006403,
  0.006429,   0.006429,    0.006429,    0.006429,
  0.006417,   0.006417,    0.006417,    0.006417,
  0.006429,   0.006429,    0.006429,    0.006429,
  0.006422,   0.006422,    0.006422,    0.006422,
  0.006422,   0.006422,    0.006422,    0.006422,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.006461,   0.006461,    0.006461,    0.006461,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.006519,   0.006519,    0.006519,    0.006519,
  0.006577,   0.006577,    0.006577,    0.006577,
  0.006596,   0.006596,    0.006596,    0.006596,
  0.006616,   0.006616,    0.006616,    0.006616,
  0.006655,   0.006655,    0.006655,    0.006655,
  0.006695,   0.006695,    0.006695,    0.006695,
  0.006732,   0.006732,    0.006732,    0.006732,
  0.006758,   0.006758,    0.006758,    0.006758,
  0.006766,   0.006766,    0.006766,    0.006766,
  0.006724,   0.006724,    0.006724,    0.006724,
  0.006682,   0.006682,    0.006682,    0.006682,
  0.006661,   0.006661,    0.006661,    0.006661,
  0.006661,   0.006661,    0.006661,    0.006661,
  0.006694,   0.006694,    0.006694,    0.006694,
  0.006631,   0.006631,    0.006631,    0.006631,
  0.006472,   0.006472,    0.006472,    0.006472,
  0.006074,   0.006074,    0.006074,    0.006074,
  0.005445,   0.005445,    0.005445,    0.005445,
  0.004988,   0.004988,    0.004988,    0.004988,
  0.004887,   0.004887,    0.004887,    0.004887,
  0.004762,   0.004762,    0.004762,    0.004762,
  0.004418,   0.004418,    0.004418,    0.004418,
  0.004177,   0.004177,    0.004177,    0.004177,
  0.004082,   0.004082,    0.004082,    0.004082,
  0.003894,   0.003894,    0.003894,    0.003894,
  0.003753,   0.003753,    0.003753,    0.003753,
  0.00369,    0.00369,     0.00369,     0.00369,
  0.003597,   0.003597,    0.003597,    0.003597,
  0.003616,   0.003616,    0.003616,    0.003616,
  0.003688,   0.003688,    0.003688,    0.003688,
  0.003746,   0.003746,    0.003746,    0.003746,
  0.003773,   0.003773,    0.003773,    0.003773,
  0.003783,   0.003783,    0.003783,    0.003783,
  0.003791,   0.003791,    0.003791,    0.003791,
  0.003809,   0.003809,    0.003809,    0.003809,
  0.003898,   0.003898,    0.003898,    0.003898,
  0.003902,   0.003902,    0.003902,    0.003902,
  0.003659,   0.003659,    0.003659,    0.003659,
  0.003382,   0.003382,    0.003382,    0.003382,
  0.003235,   0.003235,    0.003235,    0.003235,
  0.003197,   0.003197,    0.003197,    0.003197,
  0.003208,   0.003208,    0.003208,    0.003208,
  0.003224,   0.003224,    0.003224,    0.003224,
  0.003162,   0.003162,    0.003162,    0.003162,
  0.003034,   0.003034,    0.003034,    0.003034,
  0.003026,   0.003026,    0.003026,    0.003026,
  0.003096,   0.003096,    0.003096,    0.003096,
  0.003222,   0.003222,    0.003222,    0.003222,
  0.00336,    0.00336,     0.00336,     0.00336,
  0.003316,   0.003316,    0.003316,    0.003316,
  0.003285,   0.003285,    0.003285,    0.003285,
  0.003329,   0.003329,    0.003329,    0.003329,
  0.00331,    0.00331,     0.00331,     0.00331,
  0.003273,   0.003273,    0.003273,    0.003273,
  0.003204,   0.003204,    0.003204,    0.003204,
  0.003175,   0.003175,    0.003175,    0.003175,
  0.003287,   0.003287,    0.003287,    0.003287,
  0.003326,   0.003326,    0.003326,    0.003326,
  0.003272,   0.003272,    0.003272,    0.003272,
  0.003313,   0.003313,    0.003313,    0.003313,
  0.003391,   0.003391,    0.003391,    0.003391,
  0.003418,   0.003418,    0.003418,    0.003418,
  0.003389,   0.003389,    0.003389,    0.003389,
  0.003329,   0.003329,    0.003329,    0.003329,
  0.003296,   0.003296,    0.003296,    0.003296,
  0.003297,   0.003297,    0.003297,    0.003297,
  0.003236,   0.003236,    0.003236,    0.003236,
  0.003171,   0.003171,    0.003171,    0.003171,
  0.003153,   0.003153,    0.003153,    0.003153,
  0.003122,   0.003122,    0.003122,    0.003122,
  0.003187,   0.003187,    0.003187,    0.003187,
  0.003256,   0.003256,    0.003256,    0.003256,
  0.003252,   0.003252,    0.003252,    0.003252,
  0.00324,    0.00324,     0.00324,     0.00324,
  0.0032,     0.0032,      0.0032,      0.0032,
  0.003098,   0.003098,    0.003098,    0.003098,
  0.003046,   0.003046,    0.003046,    0.003046,
  0.002991,   0.002991,    0.002991,    0.002991,
  0.002945,   0.002945,    0.002945,    0.002945,
  0.002987,   0.002987,    0.002987,    0.002987,
  0.003034,   0.003034,    0.003034,    0.003034,
  0.00305,    0.00305,     0.00305,     0.00305,
  0.003024,   0.003024,    0.003024,    0.003024,
  0.003128,   0.003128,    0.003128,    0.003128,
  0.00322,    0.00322,     0.00322,     0.00322,
  0.003089,   0.003089,    0.003089,    0.003089,
  0.002769,   0.002769,    0.002769,    0.002769,
  0.002525,   0.002525,    0.002525,    0.002525,
  0.002366,   0.002366,    0.002366,    0.002366,
  0.002134,   0.002134,    0.002134,    0.002134,
  0.002036,   0.002036,    0.002036,    0.002036,
  0.002031,   0.002031,    0.002031,    0.002031,
  0.001889,   0.001889,    0.001889,    0.001889,
  0.001758,   0.001758,    0.001758,    0.001758,
  0.001735,   0.001735,    0.001735,    0.001735,
  0.001766,   0.001766,    0.001766,    0.001766,
  0.001799,   0.001799,    0.001799,    0.001799,
  0.001777,   0.001777,    0.001777,    0.001777,
  0.001801,   0.001801,    0.001801,    0.001801,
  0.001829,   0.001829,    0.001829,    0.001829,
  0.001838,   0.001838,    0.001838,    0.001838,
  0.001932,   0.001932,    0.001932,    0.001932,
  0.002018,   0.002018,    0.002018,    0.002018,
  0.002041,   0.002041,    0.002041,    0.002041,
  0.002151,   0.002151,    0.002151,    0.002151,
  0.00231,    0.00231,     0.00231,     0.00231,
  0.002416,   0.002416,    0.002416,    0.002416,
  0.002537,   0.002537,    0.002537,    0.002537,
  0.002631,   0.002631,    0.002631,    0.002631,
  0.002706,   0.002706,    0.002706,    0.002706,
  0.002698,   0.002698,    0.002698,    0.002698,
  0.002618,   0.002618,    0.002618,    0.002618,
  0.002607,   0.002607,    0.002607,    0.002607,
  0.002595,   0.002595,    0.002595,    0.002595,
  0.002581,   0.002581,    0.002581,    0.002581,
  0.002566,   0.002566,    0.002566,    0.002566,
  0.002573,   0.002573,    0.002573,    0.002573,
  0.002621,   0.002621,    0.002621,    0.002621,
  0.002628,   0.002628,    0.002628,    0.002628,
  0.002646,   0.002646,    0.002646,    0.002646,
  0.002703,   0.002703,    0.002703,    0.002703,
  0.002689,   0.002689,    0.002689,    0.002689,
  0.002653,   0.002653,    0.002653,    0.002653,
  0.002662,   0.002662,    0.002662,    0.002662,
  0.002675,   0.002675,    0.002675,    0.002675,
  0.002722,   0.002722,    0.002722,    0.002722,
  0.002757,   0.002757,    0.002757,    0.002757,
  0.002749,   0.002749,    0.002749,    0.002749,
  0.002768,   0.002768,    0.002768,    0.002768,
  0.002819,   0.002819,    0.002819,    0.002819,
  0.002811,   0.002811,    0.002811,    0.002811,
  0.002768,   0.002768,    0.002768,    0.002768,
  0.00267,    0.00267,     0.00267,     0.00267,
  0.002356,   0.002356,    0.002356,    0.002356,
  0.002091,   0.002091,    0.002091,    0.002091,
  0.001951,   0.001951,    0.001951,    0.001951,
  0.001774,   0.001774,    0.001774,    0.001774,
  0.00173,    0.00173,     0.00173,     0.00173,
  0.001729,   0.001729,    0.001729,    0.001729,
  0.00165,    0.00165,     0.00165,     0.00165,
  0.001607,   0.001607,    0.001607,    0.001607,
  0.001574,   0.001574,    0.001574,    0.001574,
  0.001452,   0.001452,    0.001452,    0.001452,
  0.00135,    0.00135,     0.00135,     0.00135,
  0.001332,   0.001332,    0.001332,    0.001332,
  0.001396,   0.001396,    0.001396,    0.001396,
  0.001547,   0.001547,    0.001547,    0.001547,
  0.001617,   0.001617,    0.001617,    0.001617,
  0.001654,   0.001654,    0.001654,    0.001654,
  0.001754,   0.001754,    0.001754,    0.001754,
  0.001825,   0.001825,    0.001825,    0.001825,
  0.001915,   0.001915,    0.001915,    0.001915,
  0.002029,   0.002029,    0.002029,    0.002029,
  0.0021,     0.0021,      0.0021,      0.0021,
  0.002197,   0.002197,    0.002197,    0.002197,
  0.002319,   0.002319,    0.002319,    0.002319,
  0.002455,   0.002455,    0.002455,    0.002455,
  0.002605,   0.002605,    0.002605,    0.002605,
  0.002706,   0.002706,    0.002706,    0.002706,
  0.002743,   0.002743,    0.002743,    0.002743,
  0.00274,    0.00274,     0.00274,     0.00274,
  0.002689,   0.002689,    0.002689,    0.002689,
  0.002645,   0.002645,    0.002645,    0.002645,
  0.002626,   0.002626,    0.002626,    0.002626,
  0.002569,   0.002569,    0.002569,    0.002569,
  0.002511,   0.002511,    0.002511,    0.002511,
  0.002493,   0.002493,    0.002493,    0.002493,
  0.002509,   0.002509,    0.002509,    0.002509,
  0.002568,   0.002568,    0.002568,    0.002568,
  0.00263,    0.00263,     0.00263,     0.00263,
  0.00267,    0.00267,     0.00267,     0.00267,
  0.002682,   0.002682,    0.002682,    0.002682,
  0.002694,   0.002694,    0.002694,    0.002694,
  0.002723,   0.002723,    0.002723,    0.002723,
  0.002768,   0.002768,    0.002768,    0.002768,
  0.002812,   0.002812,    0.002812,    0.002812,
  0.002809,   0.002809,    0.002809,    0.002809,
  0.00281,    0.00281,     0.00281,     0.00281,
  0.002846,   0.002846,    0.002846,    0.002846,
  0.002906,   0.002906,    0.002906,    0.002906,
  0.00297,    0.00297,     0.00297,     0.00297,
  0.002884,   0.002884,    0.002884,    0.002884,
  0.002779,   0.002779,    0.002779,    0.002779,
  0.002841,   0.002841,    0.002841,    0.002841,
  0.00285,    0.00285,     0.00285,     0.00285,
  0.002692,   0.002692,    0.002692,    0.002692,
  0.002387,   0.002387,    0.002387,    0.002387,
  0.002132,   0.002132,    0.002132,    0.002132,
  0.002031,   0.002031,    0.002031,    0.002031,
  0.001896,   0.001896,    0.001896,    0.001896,
  0.001667,   0.001667,    0.001667,    0.001667,
  0.001486,   0.001486,    0.001486,    0.001486,
  0.001283,   0.001283,    0.001283,    0.001283,
  0.001297,   0.001297,    0.001297,    0.001297,
  0.001626,   0.001626,    0.001626,    0.001626,
  0.001878,   0.001878,    0.001878,    0.001878,
  0.002065,   0.002065,    0.002065,    0.002065,
  0.002181,   0.002181,    0.002181,    0.002181,
  0.002238,   0.002238,    0.002238,    0.002238,
  0.002243,   0.002243,    0.002243,    0.002243,
  0.002291,   0.002291,    0.002291,    0.002291,
  0.002553,   0.002553,    0.002553,    0.002553,
  0.00307,    0.00307,     0.00307,     0.00307,
  0.003591,   0.003591,    0.003591,    0.003591,
  0.003889,   0.003889,    0.003889,    0.003889,
  0.004071,   0.004071,    0.004071,    0.004071,
  0.004206,   0.004206,    0.004206,    0.004206,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.004077,   0.004077,    0.004077,    0.004077,
  0.004186,   0.004186,    0.004186,    0.004186,
  0.004377,   0.004377,    0.004377,    0.004377,
  0.004623,   0.004623,    0.004623,    0.004623,
  0.004809,   0.004809,    0.004809,    0.004809,
  0.004902,   0.004902,    0.004902,    0.004902,
  0.004933,   0.004933,    0.004933,    0.004933,
  0.004918,   0.004918,    0.004918,    0.004918,
  0.004858,   0.004858,    0.004858,    0.004858,
  0.004696,   0.004696,    0.004696,    0.004696,
  0.004554,   0.004554,    0.004554,    0.004554,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004487,   0.004487,    0.004487,    0.004487,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004447,   0.004447,    0.004447,    0.004447,
  0.004791,   0.004791,    0.004791,    0.004791,
  0.005254,   0.005254,    0.005254,    0.005254,
  0.005686,   0.005686,    0.005686,    0.005686,
  0.005861,   0.005861,    0.005861,    0.005861,
  0.005883,   0.005883,    0.005883,    0.005883,
  0.005815,   0.005815,    0.005815,    0.005815,
  0.005605,   0.005605,    0.005605,    0.005605,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.00501,    0.00501,     0.00501,     0.00501,
  0.004968,   0.004968,    0.004968,    0.004968,
  0.004839,   0.004839,    0.004839,    0.004839,
  0.004759,   0.004759,    0.004759,    0.004759,
  0.004694,   0.004694,    0.004694,    0.004694,
  0.004739,   0.004739,    0.004739,    0.004739,
  0.004884,   0.004884,    0.004884,    0.004884,
  0.004935,   0.004935,    0.004935,    0.004935,
  0.004872,   0.004872,    0.004872,    0.004872,
  0.00469,    0.00469,     0.00469,     0.00469,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004713,   0.004713,    0.004713,    0.004713,
  0.004796,   0.004796,    0.004796,    0.004796,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004645,   0.004645,    0.004645,    0.004645,
  0.004469,   0.004469,    0.004469,    0.004469,
  0.004332,   0.004332,    0.004332,    0.004332,
  0.003985,   0.003985,    0.003985,    0.003985,
  0.003764,   0.003764,    0.003764,    0.003764,
  0.003823,   0.003823,    0.003823,    0.003823,
  0.003842,   0.003842,    0.003842,    0.003842,
  0.00391,    0.00391,     0.00391,     0.00391,
  0.004091,   0.004091,    0.004091,    0.004091,
  0.004316,   0.004316,    0.004316,    0.004316,
  0.004513,   0.004513,    0.004513,    0.004513,
  0.00465,    0.00465,     0.00465,     0.00465,
  0.00476,    0.00476,     0.00476,     0.00476,
  0.004917,   0.004917,    0.004917,    0.004917,
  0.005027,   0.005027,    0.005027,    0.005027,
  0.005059,   0.005059,    0.005059,    0.005059,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005171,   0.005171,    0.005171,    0.005171,
  0.005258,   0.005258,    0.005258,    0.005258,
  0.005333,   0.005333,    0.005333,    0.005333,
  0.005391,   0.005391,    0.005391,    0.005391,
  0.005448,   0.005448,    0.005448,    0.005448,
  0.005587,   0.005587,    0.005587,    0.005587,
  0.005751,   0.005751,    0.005751,    0.005751,
  0.005748,   0.005748,    0.005748,    0.005748,
  0.00555,    0.00555,     0.00555,     0.00555,
  0.005263,   0.005263,    0.005263,    0.005263,
  0.005082,   0.005082,    0.005082,    0.005082,
  0.005137,   0.005137,    0.005137,    0.005137,
  0.005271,   0.005271,    0.005271,    0.005271,
  0.005239,   0.005239,    0.005239,    0.005239,
  0.004991,   0.004991,    0.004991,    0.004991,
  0.004484,   0.004484,    0.004484,    0.004484,
  0.00384,    0.00384,     0.00384,     0.00384,
  0.003255,   0.003255,    0.003255,    0.003255,
  0.003035,   0.003035,    0.003035,    0.003035,
  0.003102,   0.003102,    0.003102,    0.003102,
  0.003175,   0.003175,    0.003175,    0.003175,
  0.003143,   0.003143,    0.003143,    0.003143,
  0.002941,   0.002941,    0.002941,    0.002941,
  0.002986,   0.002986,    0.002986,    0.002986,
  0.003273,   0.003273,    0.003273,    0.003273,
  0.003471,   0.003471,    0.003471,    0.003471,
  0.003579,   0.003579,    0.003579,    0.003579,
  0.003674,   0.003674,    0.003674,    0.003674,
  0.003764,   0.003764,    0.003764,    0.003764,
  0.003855,   0.003855,    0.003855,    0.003855,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003953,   0.003953,    0.003953,    0.003953,
  0.003976,   0.003976,    0.003976,    0.003976,
  0.004082,   0.004082,    0.004082,    0.004082,
  0.004128,   0.004128,    0.004128,    0.004128,
  0.004078,   0.004078,    0.004078,    0.004078,
  0.004041,   0.004041,    0.004041,    0.004041,
  0.004069,   0.004069,    0.004069,    0.004069,
  0.004069,   0.004069,    0.004069,    0.004069,
  0.004071,   0.004071,    0.004071,    0.004071,
  0.004087,   0.004087,    0.004087,    0.004087,
  0.004101,   0.004101,    0.004101,    0.004101,
  0.004054,   0.004054,    0.004054,    0.004054,
  0.00407,    0.00407,     0.00407,     0.00407,
  0.004257,   0.004257,    0.004257,    0.004257,
  0.00435,    0.00435,     0.00435,     0.00435,
  0.004461,   0.004461,    0.004461,    0.004461,
  0.004573,   0.004573,    0.004573,    0.004573,
  0.004529,   0.004529,    0.004529,    0.004529,
  0.004419,   0.004419,    0.004419,    0.004419,
  0.004354,   0.004354,    0.004354,    0.004354,
  0.004479,   0.004479,    0.004479,    0.004479,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004477,   0.004477,    0.004477,    0.004477,
  0.004341,   0.004341,    0.004341,    0.004341,
  0.00425,    0.00425,     0.00425,     0.00425,
  0.00425,    0.00425,     0.00425,     0.00425,
  0.004328,   0.004328,    0.004328,    0.004328,
  0.004345,   0.004345,    0.004345,    0.004345,
  0.004277,   0.004277,    0.004277,    0.004277,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.004326,   0.004326,    0.004326,    0.004326,
  0.003929,   0.003929,    0.003929,    0.003929,
  0.003929,   0.003929,    0.003929,    0.003929,
  0.003789,   0.003789,    0.003789,    0.003789,
  0.003587,   0.003587,    0.003587,    0.003587,
  0.0035,     0.0035,      0.0035,      0.0035,
  0.003474,   0.003474,    0.003474,    0.003474,
  0.003618,   0.003618,    0.003618,    0.003618,
  0.003744,   0.003744,    0.003744,    0.003744,
  0.003683,   0.003683,    0.003683,    0.003683,
  0.003603,   0.003603,    0.003603,    0.003603,
  0.003715,   0.003715,    0.003715,    0.003715,
  0.003981,   0.003981,    0.003981,    0.003981,
  0.004131,   0.004131,    0.004131,    0.004131,
  0.004093,   0.004093,    0.004093,    0.004093,
  0.004176,   0.004176,    0.004176,    0.004176,
  0.004495,   0.004495,    0.004495,    0.004495,
  0.004681,   0.004681,    0.004681,    0.004681,
  0.004602,   0.004602,    0.004602,    0.004602,
  0.004461,   0.004461,    0.004461,    0.004461,
  0.004384,   0.004384,    0.004384,    0.004384,
  0.004358,   0.004358,    0.004358,    0.004358,
  0.004317,   0.004317,    0.004317,    0.004317,
  0.004262,   0.004262,    0.004262,    0.004262,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004211,   0.004211,    0.004211,    0.004211,
  0.004125,   0.004125,    0.004125,    0.004125,
  0.003986,   0.003986,    0.003986,    0.003986,
  0.003877,   0.003877,    0.003877,    0.003877,
  0.003859,   0.003859,    0.003859,    0.003859,
  0.003846,   0.003846,    0.003846,    0.003846,
  0.003809,   0.003809,    0.003809,    0.003809,
  0.003853,   0.003853,    0.003853,    0.003853,
  0.003915,   0.003915,    0.003915,    0.003915,
  0.003952,   0.003952,    0.003952,    0.003952,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.003861,   0.003861,    0.003861,    0.003861,
  0.003729,   0.003729,    0.003729,    0.003729,
  0.003705,   0.003705,    0.003705,    0.003705,
  0.003788,   0.003788,    0.003788,    0.003788,
  0.003974,   0.003974,    0.003974,    0.003974,
  0.004303,   0.004303,    0.004303,    0.004303,
  0.004456,   0.004456,    0.004456,    0.004456,
  0.004345,   0.004345,    0.004345,    0.004345,
  0.004174,   0.004174,    0.004174,    0.004174,
  0.004058,   0.004058,    0.004058,    0.004058,
  0.004057,   0.004057,    0.004057,    0.004057,
  0.004025,   0.004025,    0.004025,    0.004025,
  0.003942,   0.003942,    0.003942,    0.003942,
  0.003795,   0.003795,    0.003795,    0.003795,
  0.00366,    0.00366,     0.00366,     0.00366,
  0.003731,   0.003731,    0.003731,    0.003731,
  0.003809,   0.003809,    0.003809,    0.003809,
  0.003817,   0.003817,    0.003817,    0.003817,
  0.0039,     0.0039,      0.0039,      0.0039,
  0.004057,   0.004057,    0.004057,    0.004057,
  0.004152,   0.004152,    0.004152,    0.004152,
  0.004259,   0.004259,    0.004259,    0.004259,
  0.004425,   0.004425,    0.004425,    0.004425,
  0.004498,   0.004498,    0.004498,    0.004498,
  0.00452,    0.00452,     0.00452,     0.00452,
  0.004526,   0.004526,    0.004526,    0.004526,
  0.00454,    0.00454,     0.00454,     0.00454,
  0.004593,   0.004593,    0.004593,    0.004593,
  0.004601,   0.004601,    0.004601,    0.004601,
  0.004547,   0.004547,    0.004547,    0.004547,
  0.004538,   0.004538,    0.004538,    0.004538,
  0.004611,   0.004611,    0.004611,    0.004611,
  0.00467,    0.00467,     0.00467,     0.00467,
  0.004684,   0.004684,    0.004684,    0.004684,
  0.004698,   0.004698,    0.004698,    0.004698,
  0.004726,   0.004726,    0.004726,    0.004726,
  0.004786,   0.004786,    0.004786,    0.004786,
  0.004878,   0.004878,    0.004878,    0.004878,
  0.004906,   0.004906,    0.004906,    0.004906,
  0.004921,   0.004921,    0.004921,    0.004921,
  0.004984,   0.004984,    0.004984,    0.004984,
  0.005064,   0.005064,    0.005064,    0.005064,
  0.005193,   0.005193,    0.005193,    0.005193,
  0.005339,   0.005339,    0.005339,    0.005339,
  0.005486,   0.005486,    0.005486,    0.005486,
  0.005531,   0.005531,    0.005531,    0.005531,
  0.005511,   0.005511,    0.005511,    0.005511,
  0.005508,   0.005508,    0.005508,    0.005508,
  0.005522,   0.005522,    0.005522,    0.005522,
  0.005571,   0.005571,    0.005571,    0.005571,
  0.005556,   0.005556,    0.005556,    0.005556,
  0.005595,   0.005595,    0.005595,    0.005595,
  0.005709,   0.005709,    0.005709,    0.005709,
  0.005727,   0.005727,    0.005727,    0.005727,
  0.005693,   0.005693,    0.005693,    0.005693,
  0.005629,   0.005629,    0.005629,    0.005629,
  0.005552,   0.005552,    0.005552,    0.005552,
  0.005488,   0.005488,    0.005488,    0.005488,
  0.00545,    0.00545,     0.00545,     0.00545,
  0.005423,   0.005423,    0.005423,    0.005423,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005973,   0.005973,    0.005973,    0.005973,
  0.006253,   0.006253,    0.006253,    0.006253,
  0.006246,   0.006246,    0.006246,    0.006246,
  0.00615,    0.00615,     0.00615,     0.00615,
  0.005874,   0.005874,    0.005874,    0.005874,
  0.005657,   0.005657,    0.005657,    0.005657,
  0.005495,   0.005495,    0.005495,    0.005495,
  0.005435,   0.005435,    0.005435,    0.005435,
  0.005502,   0.005502,    0.005502,    0.005502,
  0.005608,   0.005608,    0.005608,    0.005608,
  0.005565,   0.005565,    0.005565,    0.005565,
  0.005305,   0.005305,    0.005305,    0.005305,
  0.005,      0.005,       0.005,       0.005,
  0.004766,   0.004766,    0.004766,    0.004766,
  0.004719,   0.004719,    0.004719,    0.004719,
  0.004647,   0.004647,    0.004647,    0.004647,
  0.004474,   0.004474,    0.004474,    0.004474,
  0.004328,   0.004328,    0.004328,    0.004328,
  0.004122,   0.004122,    0.004122,    0.004122,
  0.003993,   0.003993,    0.003993,    0.003993,
  0.004005,   0.004005,    0.004005,    0.004005,
  0.003954,   0.003954,    0.003954,    0.003954,
  0.003854,   0.003854,    0.003854,    0.003854,
  0.003788,   0.003788,    0.003788,    0.003788,
  0.00371,    0.00371,     0.00371,     0.00371,
  0.003584,   0.003584,    0.003584,    0.003584,
  0.003441,   0.003441,    0.003441,    0.003441,
  0.003362,   0.003362,    0.003362,    0.003362,
  0.003409,   0.003409,    0.003409,    0.003409,
  0.003534,   0.003534,    0.003534,    0.003534,
  0.003658,   0.003658,    0.003658,    0.003658,
  0.003752,   0.003752,    0.003752,    0.003752,
  0.00383,    0.00383,     0.00383,     0.00383,
  0.003878,   0.003878,    0.003878,    0.003878,
  0.003816,   0.003816,    0.003816,    0.003816,
  0.003739,   0.003739,    0.003739,    0.003739,
  0.003881,   0.003881,    0.003881,    0.003881,
  0.004118,   0.004118,    0.004118,    0.004118,
  0.00418,    0.00418,     0.00418,     0.00418,
  0.004146,   0.004146,    0.004146,    0.004146,
  0.004072,   0.004072,    0.004072,    0.004072,
  0.003986,   0.003986,    0.003986,    0.003986,
  0.003933,   0.003933,    0.003933,    0.003933,
  0.003708,   0.003708,    0.003708,    0.003708,
  0.003508,   0.003508,    0.003508,    0.003508,
  0.003346,   0.003346,    0.003346,    0.003346,
  0.003251,   0.003251,    0.003251,    0.003251,
  0.00323,    0.00323,     0.00323,     0.00323,
  0.003223,   0.003223,    0.003223,    0.003223,
  0.003341,   0.003341,    0.003341,    0.003341,
  0.003329,   0.003329,    0.003329,    0.003329,
  0.003374,   0.003374,    0.003374,    0.003374,
  0.003461,   0.003461,    0.003461,    0.003461,
  0.003379,   0.003379,    0.003379,    0.003379,
  0.003278,   0.003278,    0.003278,    0.003278,
  0.003171,   0.003171,    0.003171,    0.003171,
  0.003102,   0.003102,    0.003102,    0.003102,
  0.0031,     0.0031,      0.0031,      0.0031,
  0.003206,   0.003206,    0.003206,    0.003206,
  0.003404,   0.003404,    0.003404,    0.003404,
  0.003505,   0.003505,    0.003505,    0.003505,
  0.003561,   0.003561,    0.003561,    0.003561,
  0.003475,   0.003475,    0.003475,    0.003475,
  0.003336,   0.003336,    0.003336,    0.003336,
  0.003375,   0.003375,    0.003375,    0.003375,
  0.003453,   0.003453,    0.003453,    0.003453,
  0.0035,     0.0035,      0.0035,      0.0035,
  0.003597,   0.003597,    0.003597,    0.003597,
  0.003726,   0.003726,    0.003726,    0.003726,
  0.003839,   0.003839,    0.003839,    0.003839,
  0.003952,   0.003952,    0.003952,    0.003952,
  0.004004,   0.004004,    0.004004,    0.004004,
  0.004021,   0.004021,    0.004021,    0.004021,
  0.00407,    0.00407,     0.00407,     0.00407,
  0.004155,   0.004155,    0.004155,    0.004155,
  0.004284,   0.004284,    0.004284,    0.004284,
  0.00435,    0.00435,     0.00435,     0.00435,
  0.004385,   0.004385,    0.004385,    0.004385,
  0.004427,   0.004427,    0.004427,    0.004427,
  0.004436,   0.004436,    0.004436,    0.004436,
  0.004402,   0.004402,    0.004402,    0.004402,
  0.004373,   0.004373,    0.004373,    0.004373,
  0.004402,   0.004402,    0.004402,    0.004402,
  0.004448,   0.004448,    0.004448,    0.004448,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004632,   0.004632,    0.004632,    0.004632,
  0.004706,   0.004706,    0.004706,    0.004706,
  0.004795,   0.004795,    0.004795,    0.004795,
  0.004871,   0.004871,    0.004871,    0.004871,
  0.00481,    0.00481,     0.00481,     0.00481,
  0.004627,   0.004627,    0.004627,    0.004627,
  0.004446,   0.004446,    0.004446,    0.004446,
  0.004314,   0.004314,    0.004314,    0.004314,
  0.004275,   0.004275,    0.004275,    0.004275,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004087,   0.004087,    0.004087,    0.004087,
  0.004028,   0.004028,    0.004028,    0.004028,
  0.004029,   0.004029,    0.004029,    0.004029,
  0.0039,     0.0039,      0.0039,      0.0039,
  0.004013,   0.004013,    0.004013,    0.004013,
  0.004314,   0.004314,    0.004314,    0.004314,
  0.004294,   0.004294,    0.004294,    0.004294,
  0.004207,   0.004207,    0.004207,    0.004207,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.004143,   0.004143,    0.004143,    0.004143,
  0.004143,   0.004143,    0.004143,    0.004143,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.004294,   0.004294,    0.004294,    0.004294,
  0.004356,   0.004356,    0.004356,    0.004356,
  0.004419,   0.004419,    0.004419,    0.004419,
  0.004554,   0.004554,    0.004554,    0.004554,
  0.004673,   0.004673,    0.004673,    0.004673,
  0.004818,   0.004818,    0.004818,    0.004818,
  0.004919,   0.004919,    0.004919,    0.004919,
  0.004938,   0.004938,    0.004938,    0.004938,
  0.004929,   0.004929,    0.004929,    0.004929,
  0.004844,   0.004844,    0.004844,    0.004844,
  0.00473,    0.00473,     0.00473,     0.00473,
  0.00465,    0.00465,     0.00465,     0.00465,
  0.004559,   0.004559,    0.004559,    0.004559,
  0.004471,   0.004471,    0.004471,    0.004471,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004347,   0.004347,    0.004347,    0.004347,
  0.004266,   0.004266,    0.004266,    0.004266,
  0.004187,   0.004187,    0.004187,    0.004187,
  0.004101,   0.004101,    0.004101,    0.004101,
  0.004025,   0.004025,    0.004025,    0.004025,
  0.003967,   0.003967,    0.003967,    0.003967,
  0.003932,   0.003932,    0.003932,    0.003932,
  0.003904,   0.003904,    0.003904,    0.003904,
  0.003877,   0.003877,    0.003877,    0.003877,
  0.003877,   0.003877,    0.003877,    0.003877,
  0.003908,   0.003908,    0.003908,    0.003908,
  0.00399,    0.00399,     0.00399,     0.00399,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.004312,   0.004312,    0.004312,    0.004312,
  0.004407,   0.004407,    0.004407,    0.004407,
  0.004144,   0.004144,    0.004144,    0.004144,
  0.00336,    0.00336,     0.00336,     0.00336,
  0.002386,   0.002386,    0.002386,    0.002386,
  0.001959,   0.001959,    0.001959,    0.001959,
  0.002108,   0.002108,    0.002108,    0.002108,
  0.002157,   0.002157,    0.002157,    0.002157,
  0.002042,   0.002042,    0.002042,    0.002042,
  0.002076,   0.002076,    0.002076,    0.002076,
  0.002072,   0.002072,    0.002072,    0.002072,
  0.002116,   0.002116,    0.002116,    0.002116,
  0.002258,   0.002258,    0.002258,    0.002258,
  0.002319,   0.002319,    0.002319,    0.002319,
  0.002358,   0.002358,    0.002358,    0.002358,
  0.002483,   0.002483,    0.002483,    0.002483,
  0.002657,   0.002657,    0.002657,    0.002657,
  0.002814,   0.002814,    0.002814,    0.002814,
  0.002925,   0.002925,    0.002925,    0.002925,
  0.003085,   0.003085,    0.003085,    0.003085,
  0.003237,   0.003237,    0.003237,    0.003237,
  0.003329,   0.003329,    0.003329,    0.003329,
  0.00345,    0.00345,     0.00345,     0.00345,
  0.003461,   0.003461,    0.003461,    0.003461,
  0.003421,   0.003421,    0.003421,    0.003421,
  0.003513,   0.003513,    0.003513,    0.003513,
  0.003783,   0.003783,    0.003783,    0.003783,
  0.004101,   0.004101,    0.004101,    0.004101,
  0.00427,    0.00427,     0.00427,     0.00427,
  0.004291,   0.004291,    0.004291,    0.004291,
  0.004209,   0.004209,    0.004209,    0.004209,
  0.004099,   0.004099,    0.004099,    0.004099,
  0.00401,    0.00401,     0.00401,     0.00401,
  0.003988,   0.003988,    0.003988,    0.003988,
  0.004012,   0.004012,    0.004012,    0.004012,
  0.004056,   0.004056,    0.004056,    0.004056,
  0.004134,   0.004134,    0.004134,    0.004134,
  0.004178,   0.004178,    0.004178,    0.004178,
  0.004148,   0.004148,    0.004148,    0.004148,
  0.004144,   0.004144,    0.004144,    0.004144,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004048,   0.004048,    0.004048,    0.004048,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.003752,   0.003752,    0.003752,    0.003752,
  0.003849,   0.003849,    0.003849,    0.003849,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.00401,    0.00401,     0.00401,     0.00401,
  0.004312,   0.004312,    0.004312,    0.004312,
  0.004749,   0.004749,    0.004749,    0.004749,
  0.005172,   0.005172,    0.005172,    0.005172,
  0.005352,   0.005352,    0.005352,    0.005352,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005371,   0.005371,    0.005371,    0.005371,
  0.005346,   0.005346,    0.005346,    0.005346,
  0.005325,   0.005325,    0.005325,    0.005325,
  0.005288,   0.005288,    0.005288,    0.005288,
  0.005123,   0.005123,    0.005123,    0.005123,
  0.004944,   0.004944,    0.004944,    0.004944,
  0.0049,     0.0049,      0.0049,      0.0049,
  0.004994,   0.004994,    0.004994,    0.004994,
  0.004975,   0.004975,    0.004975,    0.004975,
  0.004719,   0.004719,    0.004719,    0.004719,
  0.004513,   0.004513,    0.004513,    0.004513,
  0.004339,   0.004339,    0.004339,    0.004339,
  0.004155,   0.004155,    0.004155,    0.004155,
  0.004113,   0.004113,    0.004113,    0.004113,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004178,   0.004178,    0.004178,    0.004178,
  0.004275,   0.004275,    0.004275,    0.004275,
  0.004373,   0.004373,    0.004373,    0.004373,
  0.004433,   0.004433,    0.004433,    0.004433,
  0.004387,   0.004387,    0.004387,    0.004387,
  0.004403,   0.004403,    0.004403,    0.004403,
  0.004516,   0.004516,    0.004516,    0.004516,
  0.004605,   0.004605,    0.004605,    0.004605,
  0.004683,   0.004683,    0.004683,    0.004683,
  0.004735,   0.004735,    0.004735,    0.004735,
  0.004756,   0.004756,    0.004756,    0.004756,
  0.00471,    0.00471,     0.00471,     0.00471,
  0.004628,   0.004628,    0.004628,    0.004628,
  0.004578,   0.004578,    0.004578,    0.004578,
  0.004577,   0.004577,    0.004577,    0.004577,
  0.004575,   0.004575,    0.004575,    0.004575,
  0.004558,   0.004558,    0.004558,    0.004558,
  0.00443,    0.00443,     0.00443,     0.00443,
  0.004161,   0.004161,    0.004161,    0.004161,
  0.003957,   0.003957,    0.003957,    0.003957,
  0.0038,     0.0038,      0.0038,      0.0038,
  0.003675,   0.003675,    0.003675,    0.003675,
  0.003661,   0.003661,    0.003661,    0.003661,
  0.003661,   0.003661,    0.003661,    0.003661,
  0.003628,   0.003628,    0.003628,    0.003628,
  0.003611,   0.003611,    0.003611,    0.003611,
  0.00361,    0.00361,     0.00361,     0.00361,
  0.003579,   0.003579,    0.003579,    0.003579,
  0.003596,   0.003596,    0.003596,    0.003596,
  0.003487,   0.003487,    0.003487,    0.003487,
  0.003329,   0.003329,    0.003329,    0.003329,
  0.003266,   0.003266,    0.003266,    0.003266,
  0.003171,   0.003171,    0.003171,    0.003171,
  0.003062,   0.003062,    0.003062,    0.003062,
  0.002984,   0.002984,    0.002984,    0.002984,
  0.00297,    0.00297,     0.00297,     0.00297,
  0.002927,   0.002927,    0.002927,    0.002927,
  0.002881,   0.002881,    0.002881,    0.002881,
  0.002849,   0.002849,    0.002849,    0.002849,
  0.002881,   0.002881,    0.002881,    0.002881,
  0.002917,   0.002917,    0.002917,    0.002917,
  0.003043,   0.003043,    0.003043,    0.003043,
  0.003211,   0.003211,    0.003211,    0.003211,
  0.003141,   0.003141,    0.003141,    0.003141,
  0.003057,   0.003057,    0.003057,    0.003057,
  0.003151,   0.003151,    0.003151,    0.003151,
  0.003228,   0.003228,    0.003228,    0.003228,
  0.003159,   0.003159,    0.003159,    0.003159,
  0.00305,    0.00305,     0.00305,     0.00305,
  0.002934,   0.002934,    0.002934,    0.002934,
  0.002854,   0.002854,    0.002854,    0.002854,
  0.00292,    0.00292,     0.00292,     0.00292,
  0.003175,   0.003175,    0.003175,    0.003175,
  0.003532,   0.003532,    0.003532,    0.003532,
  0.003721,   0.003721,    0.003721,    0.003721,
  0.003847,   0.003847,    0.003847,    0.003847,
  0.003974,   0.003974,    0.003974,    0.003974,
  0.003864,   0.003864,    0.003864,    0.003864,
  0.003709,   0.003709,    0.003709,    0.003709,
  0.003686,   0.003686,    0.003686,    0.003686,
  0.003697,   0.003697,    0.003697,    0.003697,
  0.003682,   0.003682,    0.003682,    0.003682,
  0.003656,   0.003656,    0.003656,    0.003656,
  0.00363,    0.00363,     0.00363,     0.00363,
  0.003589,   0.003589,    0.003589,    0.003589,
  0.003562,   0.003562,    0.003562,    0.003562,
  0.00353,    0.00353,     0.00353,     0.00353,
  0.0035,     0.0035,      0.0035,      0.0035,
  0.003477,   0.003477,    0.003477,    0.003477,
  0.003445,   0.003445,    0.003445,    0.003445,
  0.003414,   0.003414,    0.003414,    0.003414,
  0.003408,   0.003408,    0.003408,    0.003408,
  0.003406,   0.003406,    0.003406,    0.003406,
  0.003428,   0.003428,    0.003428,    0.003428,
  0.003486,   0.003486,    0.003486,    0.003486,
  0.003527,   0.003527,    0.003527,    0.003527,
  0.00339,    0.00339,     0.00339,     0.00339,
  0.003143,   0.003143,    0.003143,    0.003143,
  0.002969,   0.002969,    0.002969,    0.002969,
  0.002697,   0.002697,    0.002697,    0.002697,
  0.002494,   0.002494,    0.002494,    0.002494,
  0.002416,   0.002416,    0.002416,    0.002416,
  0.002339,   0.002339,    0.002339,    0.002339,
  0.002174,   0.002174,    0.002174,    0.002174,
  0.001957,   0.001957,    0.001957,    0.001957,
  0.001868,   0.001868,    0.001868,    0.001868,
  0.001822,   0.001822,    0.001822,    0.001822,
  0.001757,   0.001757,    0.001757,    0.001757,
  0.00173,    0.00173,     0.00173,     0.00173,
  0.001757,   0.001757,    0.001757,    0.001757,
  0.00177,    0.00177,     0.00177,     0.00177,
  0.001798,   0.001798,    0.001798,    0.001798,
  0.001816,   0.001816,    0.001816,    0.001816,
  0.001883,   0.001883,    0.001883,    0.001883,
  0.001928,   0.001928,    0.001928,    0.001928,
  0.001938,   0.001938,    0.001938,    0.001938,
  0.001993,   0.001993,    0.001993,    0.001993,
  0.002067,   0.002067,    0.002067,    0.002067,
  0.002208,   0.002208,    0.002208,    0.002208,
  0.002354,   0.002354,    0.002354,    0.002354,
  0.002429,   0.002429,    0.002429,    0.002429,
  0.00248,    0.00248,     0.00248,     0.00248,
  0.002554,   0.002554,    0.002554,    0.002554,
  0.002647,   0.002647,    0.002647,    0.002647,
  0.002695,   0.002695,    0.002695,    0.002695,
  0.002684,   0.002684,    0.002684,    0.002684,
  0.002659,   0.002659,    0.002659,    0.002659,
  0.002631,   0.002631,    0.002631,    0.002631,
  0.00263,    0.00263,     0.00263,     0.00263,
  0.002636,   0.002636,    0.002636,    0.002636,
  0.002675,   0.002675,    0.002675,    0.002675,
  0.002733,   0.002733,    0.002733,    0.002733,
  0.002741,   0.002741,    0.002741,    0.002741,
  0.00276,    0.00276,     0.00276,     0.00276,
  0.002804,   0.002804,    0.002804,    0.002804,
  0.002811,   0.002811,    0.002811,    0.002811,
  0.002803,   0.002803,    0.002803,    0.002803,
  0.002811,   0.002811,    0.002811,    0.002811,
  0.002834,   0.002834,    0.002834,    0.002834,
  0.002834,   0.002834,    0.002834,    0.002834,
  0.002799,   0.002799,    0.002799,    0.002799,
  0.002744,   0.002744,    0.002744,    0.002744,
  0.002725,   0.002725,    0.002725,    0.002725,
  0.002749,   0.002749,    0.002749,    0.002749,
  0.002705,   0.002705,    0.002705,    0.002705,
  0.002642,   0.002642,    0.002642,    0.002642,
  0.00265,    0.00265,     0.00265,     0.00265,
  0.002656,   0.002656,    0.002656,    0.002656,
  0.002493,   0.002493,    0.002493,    0.002493,
  0.002292,   0.002292,    0.002292,    0.002292,
  0.002184,   0.002184,    0.002184,    0.002184,
  0.002099,   0.002099,    0.002099,    0.002099,
  0.002121,   0.002121,    0.002121,    0.002121,
  0.002064,   0.002064,    0.002064,    0.002064,
  0.002002,   0.002002,    0.002002,    0.002002,
  0.002041,   0.002041,    0.002041,    0.002041,
  0.002045,   0.002045,    0.002045,    0.002045,
  0.002053,   0.002053,    0.002053,    0.002053,
  0.002061,   0.002061,    0.002061,    0.002061,
  0.002153,   0.002153,    0.002153,    0.002153,
  0.002216,   0.002216,    0.002216,    0.002216,
  0.002239,   0.002239,    0.002239,    0.002239,
  0.002336,   0.002336,    0.002336,    0.002336,
  0.002584,   0.002584,    0.002584,    0.002584,
  0.002795,   0.002795,    0.002795,    0.002795,
  0.002718,   0.002718,    0.002718,    0.002718,
  0.002703,   0.002703,    0.002703,    0.002703,
  0.002908,   0.002908,    0.002908,    0.002908,
  0.00309,    0.00309,     0.00309,     0.00309,
  0.003191,   0.003191,    0.003191,    0.003191,
  0.003251,   0.003251,    0.003251,    0.003251,
  0.003298,   0.003298,    0.003298,    0.003298,
  0.003454,   0.003454,    0.003454,    0.003454,
  0.003815,   0.003815,    0.003815,    0.003815,
  0.004114,   0.004114,    0.004114,    0.004114,
  0.004178,   0.004178,    0.004178,    0.004178,
  0.004227,   0.004227,    0.004227,    0.004227,
  0.004337,   0.004337,    0.004337,    0.004337,
  0.00443,    0.00443,     0.00443,     0.00443,
  0.004429,   0.004429,    0.004429,    0.004429,
  0.004383,   0.004383,    0.004383,    0.004383,
  0.004355,   0.004355,    0.004355,    0.004355,
  0.004321,   0.004321,    0.004321,    0.004321,
  0.004291,   0.004291,    0.004291,    0.004291,
  0.00426,    0.00426,     0.00426,     0.00426,
  0.004223,   0.004223,    0.004223,    0.004223,
  0.004209,   0.004209,    0.004209,    0.004209,
  0.004196,   0.004196,    0.004196,    0.004196,
  0.004129,   0.004129,    0.004129,    0.004129,
  0.004081,   0.004081,    0.004081,    0.004081,
  0.004121,   0.004121,    0.004121,    0.004121,
  0.004241,   0.004241,    0.004241,    0.004241,
  0.004396,   0.004396,    0.004396,    0.004396,
  0.004466,   0.004466,    0.004466,    0.004466,
  0.004317,   0.004317,    0.004317,    0.004317,
  0.004035,   0.004035,    0.004035,    0.004035,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.004093,   0.004093,    0.004093,    0.004093,
  0.003696,   0.003696,    0.003696,    0.003696,
  0.003094,   0.003094,    0.003094,    0.003094,
  0.002947,   0.002947,    0.002947,    0.002947,
  0.002933,   0.002933,    0.002933,    0.002933,
  0.003041,   0.003041,    0.003041,    0.003041,
  0.003104,   0.003104,    0.003104,    0.003104,
  0.002782,   0.002782,    0.002782,    0.002782,
  0.002642,   0.002642,    0.002642,    0.002642,
  0.002781,   0.002781,    0.002781,    0.002781,
  0.002716,   0.002716,    0.002716,    0.002716,
  0.00264,    0.00264,     0.00264,     0.00264,
  0.00292,    0.00292,     0.00292,     0.00292,
  0.003185,   0.003185,    0.003185,    0.003185,
  0.003065,   0.003065,    0.003065,    0.003065,
  0.002984,   0.002984,    0.002984,    0.002984,
  0.003072,   0.003072,    0.003072,    0.003072,
  0.003193,   0.003193,    0.003193,    0.003193,
  0.003438,   0.003438,    0.003438,    0.003438,
  0.003473,   0.003473,    0.003473,    0.003473,
  0.003334,   0.003334,    0.003334,    0.003334,
  0.003328,   0.003328,    0.003328,    0.003328,
  0.003439,   0.003439,    0.003439,    0.003439,
  0.003506,   0.003506,    0.003506,    0.003506,
  0.003524,   0.003524,    0.003524,    0.003524,
  0.003528,   0.003528,    0.003528,    0.003528,
  0.003477,   0.003477,    0.003477,    0.003477,
  0.003394,   0.003394,    0.003394,    0.003394,
  0.00336,    0.00336,     0.00336,     0.00336,
  0.00333,    0.00333,     0.00333,     0.00333,
  0.003336,   0.003336,    0.003336,    0.003336,
  0.003297,   0.003297,    0.003297,    0.003297,
  0.00324,    0.00324,     0.00324,     0.00324,
  0.003384,   0.003384,    0.003384,    0.003384,
  0.003505,   0.003505,    0.003505,    0.003505,
  0.00345,    0.00345,     0.00345,     0.00345,
  0.003343,   0.003343,    0.003343,    0.003343,
  0.00326,    0.00326,     0.00326,     0.00326,
  0.00324,    0.00324,     0.00324,     0.00324,
  0.003217,   0.003217,    0.003217,    0.003217,
  0.003155,   0.003155,    0.003155,    0.003155,
  0.003141,   0.003141,    0.003141,    0.003141,
  0.003216,   0.003216,    0.003216,    0.003216,
  0.003317,   0.003317,    0.003317,    0.003317,
  0.003378,   0.003378,    0.003378,    0.003378,
  0.003377,   0.003377,    0.003377,    0.003377,
  0.003262,   0.003262,    0.003262,    0.003262,
  0.003174,   0.003174,    0.003174,    0.003174,
  0.003166,   0.003166,    0.003166,    0.003166,
  0.003072,   0.003072,    0.003072,    0.003072,
  0.002952,   0.002952,    0.002952,    0.002952,
  0.002833,   0.002833,    0.002833,    0.002833,
  0.002675,   0.002675,    0.002675,    0.002675,
  0.002587,   0.002587,    0.002587,    0.002587,
  0.002545,   0.002545,    0.002545,    0.002545,
  0.002537,   0.002537,    0.002537,    0.002537,
  0.002549,   0.002549,    0.002549,    0.002549,
  0.002447,   0.002447,    0.002447,    0.002447,
  0.002381,   0.002381,    0.002381,    0.002381,
  0.002416,   0.002416,    0.002416,    0.002416,
  0.00247,    0.00247,     0.00247,     0.00247,
  0.00253,    0.00253,     0.00253,     0.00253,
  0.002552,   0.002552,    0.002552,    0.002552,
  0.002565,   0.002565,    0.002565,    0.002565,
  0.002592,   0.002592,    0.002592,    0.002592,
  0.002554,   0.002554,    0.002554,    0.002554,
  0.002621,   0.002621,    0.002621,    0.002621,
  0.002878,   0.002878,    0.002878,    0.002878,
  0.0031,     0.0031,      0.0031,      0.0031,
  0.003204,   0.003204,    0.003204,    0.003204,
  0.003131,   0.003131,    0.003131,    0.003131,
  0.002999,   0.002999,    0.002999,    0.002999,
  0.002981,   0.002981,    0.002981,    0.002981,
  0.003014,   0.003014,    0.003014,    0.003014,
  0.002999,   0.002999,    0.002999,    0.002999,
  0.002982,   0.002982,    0.002982,    0.002982,
  0.003019,   0.003019,    0.003019,    0.003019,
  0.003107,   0.003107,    0.003107,    0.003107,
  0.003218,   0.003218,    0.003218,    0.003218,
  0.003282,   0.003282,    0.003282,    0.003282,
  0.0033,     0.0033,      0.0033,      0.0033,
  0.003287,   0.003287,    0.003287,    0.003287,
  0.003285,   0.003285,    0.003285,    0.003285,
  0.003297,   0.003297,    0.003297,    0.003297,
  0.003279,   0.003279,    0.003279,    0.003279,
  0.003264,   0.003264,    0.003264,    0.003264,
  0.003327,   0.003327,    0.003327,    0.003327,
  0.003405,   0.003405,    0.003405,    0.003405,
  0.0035,     0.0035,      0.0035,      0.0035,
  0.003648,   0.003648,    0.003648,    0.003648,
  0.003819,   0.003819,    0.003819,    0.003819,
  0.004032,   0.004032,    0.004032,    0.004032,
  0.004245,   0.004245,    0.004245,    0.004245,
  0.004395,   0.004395,    0.004395,    0.004395,
  0.004469,   0.004469,    0.004469,    0.004469,
  0.004446,   0.004446,    0.004446,    0.004446,
  0.004354,   0.004354,    0.004354,    0.004354,
  0.004287,   0.004287,    0.004287,    0.004287,
  0.004187,   0.004187,    0.004187,    0.004187,
  0.004006,   0.004006,    0.004006,    0.004006,
  0.003805,   0.003805,    0.003805,    0.003805,
  0.003607,   0.003607,    0.003607,    0.003607,
  0.003461,   0.003461,    0.003461,    0.003461,
  0.003423,   0.003423,    0.003423,    0.003423,
  0.003423,   0.003423,    0.003423,    0.003423,
  0.003311,   0.003311,    0.003311,    0.003311,
  0.003123,   0.003123,    0.003123,    0.003123,
  0.003,      0.003,       0.003,       0.003,
  0.00291,    0.00291,     0.00291,     0.00291,
  0.002874,   0.002874,    0.002874,    0.002874,
  0.002973,   0.002973,    0.002973,    0.002973,
  0.003015,   0.003015,    0.003015,    0.003015,
  0.002923,   0.002923,    0.002923,    0.002923,
  0.002973,   0.002973,    0.002973,    0.002973,
  0.003108,   0.003108,    0.003108,    0.003108,
  0.003256,   0.003256,    0.003256,    0.003256,
  0.003426,   0.003426,    0.003426,    0.003426,
  0.003557,   0.003557,    0.003557,    0.003557,
  0.00362,    0.00362,     0.00362,     0.00362,
  0.003701,   0.003701,    0.003701,    0.003701,
  0.003879,   0.003879,    0.003879,    0.003879,
  0.00405,    0.00405,     0.00405,     0.00405,
  0.0042,     0.0042,      0.0042,      0.0042,
  0.004392,   0.004392,    0.004392,    0.004392,
  0.004569,   0.004569,    0.004569,    0.004569,
  0.004697,   0.004697,    0.004697,    0.004697,
  0.004816,   0.004816,    0.004816,    0.004816,
  0.004929,   0.004929,    0.004929,    0.004929,
  0.005049,   0.005049,    0.005049,    0.005049,
  0.005149,   0.005149,    0.005149,    0.005149,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005189,   0.005189,    0.005189,    0.005189,
  0.005228,   0.005228,    0.005228,    0.005228,
  0.005231,   0.005231,    0.005231,    0.005231,
  0.005235,   0.005235,    0.005235,    0.005235,
  0.005231,   0.005231,    0.005231,    0.005231,
  0.005235,   0.005235,    0.005235,    0.005235,
  0.005312,   0.005312,    0.005312,    0.005312,
  0.005447,   0.005447,    0.005447,    0.005447,
  0.005546,   0.005546,    0.005546,    0.005546,
  0.00563,    0.00563,     0.00563,     0.00563,
  0.005751,   0.005751,    0.005751,    0.005751,
  0.005866,   0.005866,    0.005866,    0.005866,
  0.005947,   0.005947,    0.005947,    0.005947,
  0.005949,   0.005949,    0.005949,    0.005949,
  0.005858,   0.005858,    0.005858,    0.005858,
  0.00583,    0.00583,     0.00583,     0.00583,
  0.005905,   0.005905,    0.005905,    0.005905,
  0.005823,   0.005823,    0.005823,    0.005823,
  0.005859,   0.005859,    0.005859,    0.005859,
  0.006367,   0.006367,    0.006367,    0.006367,
  0.00682,    0.00682,     0.00682,     0.00682,
  0.006903,   0.006903,    0.006903,    0.006903,
  0.006924,   0.006924,    0.006924,    0.006924,
  0.006872,   0.006872,    0.006872,    0.006872,
  0.006768,   0.006768,    0.006768,    0.006768,
  0.006715,   0.006715,    0.006715,    0.006715,
  0.006693,   0.006693,    0.006693,    0.006693,
  0.006692,   0.006692,    0.006692,    0.006692,
  0.00664,    0.00664,     0.00664,     0.00664,
  0.006629,   0.006629,    0.006629,    0.006629,
  0.006641,   0.006641,    0.006641,    0.006641,
  0.006633,   0.006633,    0.006633,    0.006633,
  0.006563,   0.006563,    0.006563,    0.006563,
  0.006443,   0.006443,    0.006443,    0.006443,
  0.006364,   0.006364,    0.006364,    0.006364,
  0.006305,   0.006305,    0.006305,    0.006305,
  0.006259,   0.006259,    0.006259,    0.006259,
  0.006246,   0.006246,    0.006246,    0.006246,
  0.006214,   0.006214,    0.006214,    0.006214,
  0.006184,   0.006184,    0.006184,    0.006184,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.006104,   0.006104,    0.006104,    0.006104,
  0.006104,   0.006104,    0.006104,    0.006104,
  0.006086,   0.006086,    0.006086,    0.006086,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.005871,   0.005871,    0.005871,    0.005871,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005749,   0.005749,    0.005749,    0.005749,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005682,   0.005682,    0.005682,    0.005682,
  0.005755,   0.005755,    0.005755,    0.005755,
  0.005939,   0.005939,    0.005939,    0.005939,
  0.006058,   0.006058,    0.006058,    0.006058,
  0.006062,   0.006062,    0.006062,    0.006062,
  0.006057,   0.006057,    0.006057,    0.006057,
  0.006033,   0.006033,    0.006033,    0.006033,
  0.006039,   0.006039,    0.006039,    0.006039,
  0.005967,   0.005967,    0.005967,    0.005967,
  0.005756,   0.005756,    0.005756,    0.005756,
  0.00558,    0.00558,     0.00558,     0.00558,
  0.005476,   0.005476,    0.005476,    0.005476,
  0.005399,   0.005399,    0.005399,    0.005399,
  0.00535,    0.00535,     0.00535,     0.00535,
  0.005339,   0.005339,    0.005339,    0.005339,
  0.005377,   0.005377,    0.005377,    0.005377,
  0.005346,   0.005346,    0.005346,    0.005346,
  0.00539,    0.00539,     0.00539,     0.00539,
  0.005484,   0.005484,    0.005484,    0.005484,
  0.005354,   0.005354,    0.005354,    0.005354,
  0.005316,   0.005316,    0.005316,    0.005316,
  0.005491,   0.005491,    0.005491,    0.005491,
  0.005472,   0.005472,    0.005472,    0.005472,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005515,   0.005515,    0.005515,    0.005515,
  0.005636,   0.005636,    0.005636,    0.005636,
  0.00571,    0.00571,     0.00571,     0.00571,
  0.005721,   0.005721,    0.005721,    0.005721,
  0.005791,   0.005791,    0.005791,    0.005791,
  0.006202,   0.006202,    0.006202,    0.006202,
  0.006762,   0.006762,    0.006762,    0.006762,
  0.00705,    0.00705,     0.00705,     0.00705,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.007018,   0.007018,    0.007018,    0.007018,
  0.00705,    0.00705,     0.00705,     0.00705,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.007039,   0.007039,    0.007039,    0.007039,
  0.006998,   0.006998,    0.006998,    0.006998,
  0.006937,   0.006937,    0.006937,    0.006937,
  0.006896,   0.006896,    0.006896,    0.006896,
  0.006875,   0.006875,    0.006875,    0.006875,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006835,   0.006835,    0.006835,    0.006835,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006875,   0.006875,    0.006875,    0.006875,
  0.006875,   0.006875,    0.006875,    0.006875,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006835,   0.006835,    0.006835,    0.006835,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006875,   0.006875,    0.006875,    0.006875,
  0.006896,   0.006896,    0.006896,    0.006896,
  0.006957,   0.006957,    0.006957,    0.006957,
  0.007019,   0.007019,    0.007019,    0.007019,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.00725,    0.00725,     0.00725,     0.00725,
  0.00739,    0.00739,     0.00739,     0.00739,
  0.007444,   0.007444,    0.007444,    0.007444,
  0.007378,   0.007378,    0.007378,    0.007378,
  0.007233,   0.007233,    0.007233,    0.007233,
  0.007076,   0.007076,    0.007076,    0.007076,
  0.006994,   0.006994,    0.006994,    0.006994,
  0.007085,   0.007085,    0.007085,    0.007085,
  0.007148,   0.007148,    0.007148,    0.007148,
  0.007085,   0.007085,    0.007085,    0.007085,
  0.006946,   0.006946,    0.006946,    0.006946,
  0.00696,    0.00696,     0.00696,     0.00696,
  0.007306,   0.007306,    0.007306,    0.007306,
  0.007611,   0.007611,    0.007611,    0.007611,
  0.007698,   0.007698,    0.007698,    0.007698,
  0.007663,   0.007663,    0.007663,    0.007663,
  0.007475,   0.007475,    0.007475,    0.007475,
  0.007323,   0.007323,    0.007323,    0.007323,
  0.007305,   0.007305,    0.007305,    0.007305,
  0.007373,   0.007373,    0.007373,    0.007373,
  0.007374,   0.007374,    0.007374,    0.007374,
  0.007232,   0.007232,    0.007232,    0.007232,
  0.007167,   0.007167,    0.007167,    0.007167,
  0.007169,   0.007169,    0.007169,    0.007169,
  0.007121,   0.007121,    0.007121,    0.007121,
  0.007034,   0.007034,    0.007034,    0.007034,
  0.006946,   0.006946,    0.006946,    0.006946,
  0.006821,   0.006821,    0.006821,    0.006821,
  0.006801,   0.006801,    0.006801,    0.006801,
  0.006874,   0.006874,    0.006874,    0.006874,
  0.006915,   0.006915,    0.006915,    0.006915,
  0.006977,   0.006977,    0.006977,    0.006977,
  0.007018,   0.007018,    0.007018,    0.007018,
  0.006925,   0.006925,    0.006925,    0.006925,
  0.006831,   0.006831,    0.006831,    0.006831,
  0.006831,   0.006831,    0.006831,    0.006831,
  0.0068,     0.0068,      0.0068,      0.0068,
  0.006759,   0.006759,    0.006759,    0.006759,
  0.006709,   0.006709,    0.006709,    0.006709,
  0.006601,   0.006601,    0.006601,    0.006601,
  0.006514,   0.006514,    0.006514,    0.006514,
  0.00647,    0.00647,     0.00647,     0.00647,
  0.006455,   0.006455,    0.006455,    0.006455,
  0.006489,   0.006489,    0.006489,    0.006489,
  0.006601,   0.006601,    0.006601,    0.006601,
  0.006741,   0.006741,    0.006741,    0.006741,
  0.006835,   0.006835,    0.006835,    0.006835,
  0.006937,   0.006937,    0.006937,    0.006937,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.007186,   0.007186,    0.007186,    0.007186,
  0.007335,   0.007335,    0.007335,    0.007335,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.007597,   0.007597,    0.007597,    0.007597,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007799,   0.007799,    0.007799,    0.007799,
  0.00789,    0.00789,     0.00789,     0.00789,
  0.007904,   0.007904,    0.007904,    0.007904,
  0.007942,   0.007942,    0.007942,    0.007942,
  0.008021,   0.008021,    0.008021,    0.008021,
  0.007991,   0.007991,    0.007991,    0.007991,
  0.00789,    0.00789,     0.00789,     0.00789,
  0.007792,   0.007792,    0.007792,    0.007792,
  0.00747,    0.00747,     0.00747,     0.00747,
  0.007017,   0.007017,    0.007017,    0.007017,
  0.006808,   0.006808,    0.006808,    0.006808,
  0.006801,   0.006801,    0.006801,    0.006801,
  0.006832,   0.006832,    0.006832,    0.006832,
  0.00683,    0.00683,     0.00683,     0.00683,
  0.006766,   0.006766,    0.006766,    0.006766,
  0.006757,   0.006757,    0.006757,    0.006757,
  0.006915,   0.006915,    0.006915,    0.006915,
  0.007092,   0.007092,    0.007092,    0.007092,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007133,   0.007133,    0.007133,    0.007133,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007186,   0.007186,    0.007186,    0.007186,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007218,   0.007218,    0.007218,    0.007218,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.006997,   0.006997,    0.006997,    0.006997,
  0.006894,   0.006894,    0.006894,    0.006894,
  0.006801,   0.006801,    0.006801,    0.006801,
  0.006698,   0.006698,    0.006698,    0.006698,
  0.006583,   0.006583,    0.006583,    0.006583,
  0.0065,     0.0065,      0.0065,      0.0065,
  0.006468,   0.006468,    0.006468,    0.006468,
  0.006457,   0.006457,    0.006457,    0.006457,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.006514,   0.006514,    0.006514,    0.006514,
  0.006549,   0.006549,    0.006549,    0.006549,
  0.006584,   0.006584,    0.006584,    0.006584,
  0.006596,   0.006596,    0.006596,    0.006596,
  0.006616,   0.006616,    0.006616,    0.006616,
  0.006624,   0.006624,    0.006624,    0.006624,
  0.006632,   0.006632,    0.006632,    0.006632,
  0.006652,   0.006652,    0.006652,    0.006652,
  0.006644,   0.006644,    0.006644,    0.006644,
  0.006636,   0.006636,    0.006636,    0.006636,
  0.006624,   0.006624,    0.006624,    0.006624,
  0.006632,   0.006632,    0.006632,    0.006632,
  0.006617,   0.006617,    0.006617,    0.006617,
  0.006581,   0.006581,    0.006581,    0.006581,
  0.006537,   0.006537,    0.006537,    0.006537,
  0.006494,   0.006494,    0.006494,    0.006494,
  0.006494,   0.006494,    0.006494,    0.006494,
  0.006474,   0.006474,    0.006474,    0.006474,
  0.006444,   0.006444,    0.006444,    0.006444,
  0.006363,   0.006363,    0.006363,    0.006363,
  0.006279,   0.006279,    0.006279,    0.006279,
  0.006279,   0.006279,    0.006279,    0.006279,
  0.006329,   0.006329,    0.006329,    0.006329,
  0.006354,   0.006354,    0.006354,    0.006354,
  0.006353,   0.006353,    0.006353,    0.006353,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006327,   0.006327,    0.006327,    0.006327,
  0.006327,   0.006327,    0.006327,    0.006327,
  0.006327,   0.006327,    0.006327,    0.006327,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006384,   0.006384,    0.006384,    0.006384,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006234,   0.006234,    0.006234,    0.006234,
  0.006123,   0.006123,    0.006123,    0.006123,
  0.006014,   0.006014,    0.006014,    0.006014,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.005801,   0.005801,    0.005801,    0.005801,
  0.005748,   0.005748,    0.005748,    0.005748,
  0.005714,   0.005714,    0.005714,    0.005714,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005784,   0.005784,    0.005784,    0.005784,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006179,   0.006179,    0.006179,    0.006179,
  0.006353,   0.006353,    0.006353,    0.006353,
  0.006361,   0.006361,    0.006361,    0.006361,
  0.006218,   0.006218,    0.006218,    0.006218,
  0.006132,   0.006132,    0.006132,    0.006132,
  0.006128,   0.006128,    0.006128,    0.006128,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.006152,   0.006152,    0.006152,    0.006152,
  0.006148,   0.006148,    0.006148,    0.006148,
  0.006155,   0.006155,    0.006155,    0.006155,
  0.00621,    0.00621,     0.00621,     0.00621,
  0.006178,   0.006178,    0.006178,    0.006178,
  0.006098,   0.006098,    0.006098,    0.006098,
  0.006129,   0.006129,    0.006129,    0.006129,
  0.006153,   0.006153,    0.006153,    0.006153,
  0.006193,   0.006193,    0.006193,    0.006193,
  0.006279,   0.006279,    0.006279,    0.006279,
  0.006311,   0.006311,    0.006311,    0.006311,
  0.006284,   0.006284,    0.006284,    0.006284,
  0.006247,   0.006247,    0.006247,    0.006247,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006353,   0.006353,    0.006353,    0.006353,
  0.006312,   0.006312,    0.006312,    0.006312,
  0.006239,   0.006239,    0.006239,    0.006239,
  0.006227,   0.006227,    0.006227,    0.006227,
  0.00615,    0.00615,     0.00615,     0.00615,
  0.006157,   0.006157,    0.006157,    0.006157,
  0.006199,   0.006199,    0.006199,    0.006199,
  0.006172,   0.006172,    0.006172,    0.006172,
  0.00614,    0.00614,     0.00614,     0.00614,
  0.006097,   0.006097,    0.006097,    0.006097,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.005912,   0.005912,    0.005912,    0.005912,
  0.005835,   0.005835,    0.005835,    0.005835,
  0.005847,   0.005847,    0.005847,    0.005847,
  0.005739,   0.005739,    0.005739,    0.005739,
  0.005597,   0.005597,    0.005597,    0.005597,
  0.00556,    0.00556,     0.00556,     0.00556,
  0.005461,   0.005461,    0.005461,    0.005461,
  0.005266,   0.005266,    0.005266,    0.005266,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004759,   0.004759,    0.004759,    0.004759,
  0.004614,   0.004614,    0.004614,    0.004614,
  0.004585,   0.004585,    0.004585,    0.004585,
  0.004642,   0.004642,    0.004642,    0.004642,
  0.004896,   0.004896,    0.004896,    0.004896,
  0.005401,   0.005401,    0.005401,    0.005401,
  0.005929,   0.005929,    0.005929,    0.005929,
  0.006348,   0.006348,    0.006348,    0.006348,
  0.006677,   0.006677,    0.006677,    0.006677,
  0.007012,   0.007012,    0.007012,    0.007012,
  0.006849,   0.006849,    0.006849,    0.006849,
  0.006439,   0.006439,    0.006439,    0.006439,
  0.006275,   0.006275,    0.006275,    0.006275,
  0.006133,   0.006133,    0.006133,    0.006133,
  0.006125,   0.006125,    0.006125,    0.006125,
  0.006118,   0.006118,    0.006118,    0.006118,
  0.0061,     0.0061,      0.0061,      0.0061,
  0.006152,   0.006152,    0.006152,    0.006152,
  0.006123,   0.006123,    0.006123,    0.006123,
  0.00599,    0.00599,     0.00599,     0.00599,
  0.005751,   0.005751,    0.005751,    0.005751,
  0.005596,   0.005596,    0.005596,    0.005596,
  0.005692,   0.005692,    0.005692,    0.005692,
  0.005752,   0.005752,    0.005752,    0.005752,
  0.005687,   0.005687,    0.005687,    0.005687,
  0.005684,   0.005684,    0.005684,    0.005684,
  0.005682,   0.005682,    0.005682,    0.005682,
  0.005618,   0.005618,    0.005618,    0.005618,
  0.005745,   0.005745,    0.005745,    0.005745,
  0.006102,   0.006102,    0.006102,    0.006102,
  0.006319,   0.006319,    0.006319,    0.006319,
  0.006385,   0.006385,    0.006385,    0.006385,
  0.006484,   0.006484,    0.006484,    0.006484,
  0.006518,   0.006518,    0.006518,    0.006518,
  0.006488,   0.006488,    0.006488,    0.006488,
  0.00651,    0.00651,     0.00651,     0.00651,
  0.00657,    0.00657,     0.00657,     0.00657,
  0.006615,   0.006615,    0.006615,    0.006615,
  0.006642,   0.006642,    0.006642,    0.006642,
  0.006674,   0.006674,    0.006674,    0.006674,
  0.006683,   0.006683,    0.006683,    0.006683,
  0.006625,   0.006625,    0.006625,    0.006625,
  0.006599,   0.006599,    0.006599,    0.006599,
  0.006567,   0.006567,    0.006567,    0.006567,
  0.006493,   0.006493,    0.006493,    0.006493,
  0.006431,   0.006431,    0.006431,    0.006431,
  0.006355,   0.006355,    0.006355,    0.006355,
  0.006255,   0.006255,    0.006255,    0.006255,
  0.006121,   0.006121,    0.006121,    0.006121,
  0.006065,   0.006065,    0.006065,    0.006065,
  0.00606,    0.00606,     0.00606,     0.00606,
  0.006097,   0.006097,    0.006097,    0.006097,
  0.006292,   0.006292,    0.006292,    0.006292,
  0.006651,   0.006651,    0.006651,    0.006651,
  0.006886,   0.006886,    0.006886,    0.006886,
  0.006901,   0.006901,    0.006901,    0.006901,
  0.006819,   0.006819,    0.006819,    0.006819,
  0.006604,   0.006604,    0.006604,    0.006604,
  0.006488,   0.006488,    0.006488,    0.006488,
  0.006368,   0.006368,    0.006368,    0.006368,
  0.006128,   0.006128,    0.006128,    0.006128,
  0.0059,     0.0059,      0.0059,      0.0059,
  0.005589,   0.005589,    0.005589,    0.005589,
  0.005445,   0.005445,    0.005445,    0.005445,
  0.005317,   0.005317,    0.005317,    0.005317,
  0.005126,   0.005126,    0.005126,    0.005126,
  0.005163,   0.005163,    0.005163,    0.005163,
  0.005257,   0.005257,    0.005257,    0.005257,
  0.005204,   0.005204,    0.005204,    0.005204,
  0.005119,   0.005119,    0.005119,    0.005119,
  0.005136,   0.005136,    0.005136,    0.005136,
  0.005184,   0.005184,    0.005184,    0.005184,
  0.005246,   0.005246,    0.005246,    0.005246,
  0.005252,   0.005252,    0.005252,    0.005252,
  0.005342,   0.005342,    0.005342,    0.005342,
  0.005776,   0.005776,    0.005776,    0.005776,
  0.006258,   0.006258,    0.006258,    0.006258,
  0.006543,   0.006543,    0.006543,    0.006543,
  0.006727,   0.006727,    0.006727,    0.006727,
  0.006767,   0.006767,    0.006767,    0.006767,
  0.006713,   0.006713,    0.006713,    0.006713,
  0.006692,   0.006692,    0.006692,    0.006692,
  0.006796,   0.006796,    0.006796,    0.006796,
  0.006791,   0.006791,    0.006791,    0.006791,
  0.00677,    0.00677,     0.00677,     0.00677,
  0.006882,   0.006882,    0.006882,    0.006882,
  0.006916,   0.006916,    0.006916,    0.006916,
  0.006954,   0.006954,    0.006954,    0.006954,
  0.007007,   0.007007,    0.007007,    0.007007,
  0.006815,   0.006815,    0.006815,    0.006815,
  0.006584,   0.006584,    0.006584,    0.006584,
  0.006649,   0.006649,    0.006649,    0.006649,
  0.006673,   0.006673,    0.006673,    0.006673,
  0.00663,    0.00663,     0.00663,     0.00663,
  0.006654,   0.006654,    0.006654,    0.006654,
  0.006677,   0.006677,    0.006677,    0.006677,
  0.006669,   0.006669,    0.006669,    0.006669,
  0.006561,   0.006561,    0.006561,    0.006561,
  0.00657,    0.00657,     0.00657,     0.00657,
  0.006518,   0.006518,    0.006518,    0.006518,
  0.006442,   0.006442,    0.006442,    0.006442,
  0.006649,   0.006649,    0.006649,    0.006649,
  0.006923,   0.006923,    0.006923,    0.006923,
  0.006853,   0.006853,    0.006853,    0.006853,
  0.006583,   0.006583,    0.006583,    0.006583,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.006414,   0.006414,    0.006414,    0.006414,
  0.006433,   0.006433,    0.006433,    0.006433,
  0.006413,   0.006413,    0.006413,    0.006413,
  0.006373,   0.006373,    0.006373,    0.006373,
  0.006246,   0.006246,    0.006246,    0.006246,
  0.006063,   0.006063,    0.006063,    0.006063,
  0.005888,   0.005888,    0.005888,    0.005888,
  0.005786,   0.005786,    0.005786,    0.005786,
  0.005698,   0.005698,    0.005698,    0.005698,
  0.005571,   0.005571,    0.005571,    0.005571,
  0.00542,    0.00542,     0.00542,     0.00542,
  0.00531,    0.00531,     0.00531,     0.00531,
  0.005309,   0.005309,    0.005309,    0.005309,
  0.005417,   0.005417,    0.005417,    0.005417,
  0.005692,   0.005692,    0.005692,    0.005692,
  0.006063,   0.006063,    0.006063,    0.006063,
  0.006391,   0.006391,    0.006391,    0.006391,
  0.006536,   0.006536,    0.006536,    0.006536,
  0.006602,   0.006602,    0.006602,    0.006602,
  0.006657,   0.006657,    0.006657,    0.006657,
  0.006634,   0.006634,    0.006634,    0.006634,
  0.006653,   0.006653,    0.006653,    0.006653,
  0.006674,   0.006674,    0.006674,    0.006674,
  0.006632,   0.006632,    0.006632,    0.006632,
  0.006522,   0.006522,    0.006522,    0.006522,
  0.006352,   0.006352,    0.006352,    0.006352,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006358,   0.006358,    0.006358,    0.006358,
  0.006414,   0.006414,    0.006414,    0.006414,
  0.00647,    0.00647,     0.00647,     0.00647,
  0.006491,   0.006491,    0.006491,    0.006491,
  0.006551,   0.006551,    0.006551,    0.006551,
  0.006618,   0.006618,    0.006618,    0.006618,
  0.006674,   0.006674,    0.006674,    0.006674,
  0.006732,   0.006732,    0.006732,    0.006732,
  0.006773,   0.006773,    0.006773,    0.006773,
  0.006857,   0.006857,    0.006857,    0.006857,
  0.007008,   0.007008,    0.007008,    0.007008,
  0.007225,   0.007225,    0.007225,    0.007225,
  0.007488,   0.007488,    0.007488,    0.007488,
  0.007697,   0.007697,    0.007697,    0.007697,
  0.007799,   0.007799,    0.007799,    0.007799,
  0.007806,   0.007806,    0.007806,    0.007806,
  0.007757,   0.007757,    0.007757,    0.007757,
  0.007725,   0.007725,    0.007725,    0.007725,
  0.007715,   0.007715,    0.007715,    0.007715,
  0.007674,   0.007674,    0.007674,    0.007674,
  0.007611,   0.007611,    0.007611,    0.007611,
  0.007632,   0.007632,    0.007632,    0.007632,
  0.007707,   0.007707,    0.007707,    0.007707,
  0.007496,   0.007496,    0.007496,    0.007496,
  0.007364,   0.007364,    0.007364,    0.007364,
  0.00747,    0.00747,     0.00747,     0.00747,
  0.00742,    0.00742,     0.00742,     0.00742,
  0.007299,   0.007299,    0.007299,    0.007299,
  0.007326,   0.007326,    0.007326,    0.007326,
  0.007544,   0.007544,    0.007544,    0.007544,
  0.007635,   0.007635,    0.007635,    0.007635,
  0.007961,   0.007961,    0.007961,    0.007961,
  0.008637,   0.008637,    0.008637,    0.008637,
  0.008841,   0.008841,    0.008841,    0.008841,
  0.008956,   0.008956,    0.008956,    0.008956,
  0.009198,   0.009198,    0.009198,    0.009198,
  0.009217,   0.009217,    0.009217,    0.009217,
  0.009227,   0.009227,    0.009227,    0.009227,
  0.009205,   0.009205,    0.009205,    0.009205,
  0.0092,     0.0092,      0.0092,      0.0092,
  0.009185,   0.009185,    0.009185,    0.009185,
  0.009117,   0.009117,    0.009117,    0.009117,
  0.009077,   0.009077,    0.009077,    0.009077,
  0.009031,   0.009031,    0.009031,    0.009031,
  0.00896,    0.00896,     0.00896,     0.00896,
  0.008438,   0.008438,    0.008438,    0.008438,
  0.007605,   0.007605,    0.007605,    0.007605,
  0.007294,   0.007294,    0.007294,    0.007294,
  0.007268,   0.007268,    0.007268,    0.007268,
  0.00711,    0.00711,     0.00711,     0.00711,
  0.006989,   0.006989,    0.006989,    0.006989,
  0.006972,   0.006972,    0.006972,    0.006972,
  0.007004,   0.007004,    0.007004,    0.007004,
  0.007046,   0.007046,    0.007046,    0.007046,
  0.007092,   0.007092,    0.007092,    0.007092,
  0.007164,   0.007164,    0.007164,    0.007164,
  0.007191,   0.007191,    0.007191,    0.007191,
  0.00718,    0.00718,     0.00718,     0.00718,
  0.007226,   0.007226,    0.007226,    0.007226,
  0.007297,   0.007297,    0.007297,    0.007297,
  0.007392,   0.007392,    0.007392,    0.007392,
  0.007541,   0.007541,    0.007541,    0.007541,
  0.007642,   0.007642,    0.007642,    0.007642,
  0.007665,   0.007665,    0.007665,    0.007665,
  0.007634,   0.007634,    0.007634,    0.007634,
  0.007587,   0.007587,    0.007587,    0.007587,
  0.00766,    0.00766,     0.00766,     0.00766,
  0.0077,     0.0077,      0.0077,      0.0077,
  0.007755,   0.007755,    0.007755,    0.007755,
  0.008151,   0.008151,    0.008151,    0.008151,
  0.008395,   0.008395,    0.008395,    0.008395,
  0.008193,   0.008193,    0.008193,    0.008193,
  0.007974,   0.007974,    0.007974,    0.007974,
  0.007746,   0.007746,    0.007746,    0.007746,
  0.007536,   0.007536,    0.007536,    0.007536,
  0.007441,   0.007441,    0.007441,    0.007441,
  0.007301,   0.007301,    0.007301,    0.007301,
  0.007416,   0.007416,    0.007416,    0.007416,
  0.007534,   0.007534,    0.007534,    0.007534,
  0.00744,    0.00744,     0.00744,     0.00744,
  0.007557,   0.007557,    0.007557,    0.007557,
  0.007759,   0.007759,    0.007759,    0.007759,
  0.00788,    0.00788,     0.00788,     0.00788,
  0.007817,   0.007817,    0.007817,    0.007817,
  0.007704,   0.007704,    0.007704,    0.007704,
  0.007639,   0.007639,    0.007639,    0.007639,
  0.007594,   0.007594,    0.007594,    0.007594,
  0.007657,   0.007657,    0.007657,    0.007657,
  0.007733,   0.007733,    0.007733,    0.007733,
  0.007767,   0.007767,    0.007767,    0.007767,
  0.007762,   0.007762,    0.007762,    0.007762,
  0.00769,    0.00769,     0.00769,     0.00769,
  0.007638,   0.007638,    0.007638,    0.007638,
  0.00761,    0.00761,     0.00761,     0.00761,
  0.007569,   0.007569,    0.007569,    0.007569,
  0.007512,   0.007512,    0.007512,    0.007512,
  0.007535,   0.007535,    0.007535,    0.007535,
  0.007646,   0.007646,    0.007646,    0.007646,
  0.007681,   0.007681,    0.007681,    0.007681,
  0.007654,   0.007654,    0.007654,    0.007654,
  0.007641,   0.007641,    0.007641,    0.007641,
  0.007731,   0.007731,    0.007731,    0.007731,
  0.007867,   0.007867,    0.007867,    0.007867,
  0.007768,   0.007768,    0.007768,    0.007768,
  0.007447,   0.007447,    0.007447,    0.007447,
  0.007282,   0.007282,    0.007282,    0.007282,
  0.007357,   0.007357,    0.007357,    0.007357,
  0.007465,   0.007465,    0.007465,    0.007465,
  0.007531,   0.007531,    0.007531,    0.007531,
  0.007531,   0.007531,    0.007531,    0.007531,
  0.007172,   0.007172,    0.007172,    0.007172,
  0.006506,   0.006506,    0.006506,    0.006506,
  0.005998,   0.005998,    0.005998,    0.005998,
  0.005732,   0.005732,    0.005732,    0.005732,
  0.005578,   0.005578,    0.005578,    0.005578,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.005315,   0.005315,    0.005315,    0.005315,
  0.0053,     0.0053,      0.0053,      0.0053,
  0.005331,   0.005331,    0.005331,    0.005331,
  0.005348,   0.005348,    0.005348,    0.005348,
  0.005316,   0.005316,    0.005316,    0.005316,
  0.005219,   0.005219,    0.005219,    0.005219,
  0.00517,    0.00517,     0.00517,     0.00517,
  0.005059,   0.005059,    0.005059,    0.005059,
  0.004949,   0.004949,    0.004949,    0.004949,
  0.004949,   0.004949,    0.004949,    0.004949,
  0.004965,   0.004965,    0.004965,    0.004965,
  0.00498,    0.00498,     0.00498,     0.00498,
  0.004949,   0.004949,    0.004949,    0.004949,
  0.004886,   0.004886,    0.004886,    0.004886,
  0.004808,   0.004808,    0.004808,    0.004808,
  0.004687,   0.004687,    0.004687,    0.004687,
  0.004611,   0.004611,    0.004611,    0.004611,
  0.004284,   0.004284,    0.004284,    0.004284,
  0.003893,   0.003893,    0.003893,    0.003893,
  0.003843,   0.003843,    0.003843,    0.003843,
  0.003884,   0.003884,    0.003884,    0.003884,
  0.004006,   0.004006,    0.004006,    0.004006,
  0.004184,   0.004184,    0.004184,    0.004184,
  0.004254,   0.004254,    0.004254,    0.004254,
  0.004239,   0.004239,    0.004239,    0.004239,
  0.004164,   0.004164,    0.004164,    0.004164,
  0.004015,   0.004015,    0.004015,    0.004015,
  0.003881,   0.003881,    0.003881,    0.003881,
  0.003821,   0.003821,    0.003821,    0.003821,
  0.003825,   0.003825,    0.003825,    0.003825,
  0.003864,   0.003864,    0.003864,    0.003864,
  0.003904,   0.003904,    0.003904,    0.003904,
  0.003891,   0.003891,    0.003891,    0.003891,
  0.003879,   0.003879,    0.003879,    0.003879,
  0.003929,   0.003929,    0.003929,    0.003929,
  0.003987,   0.003987,    0.003987,    0.003987,
  0.003954,   0.003954,    0.003954,    0.003954,
  0.003839,   0.003839,    0.003839,    0.003839,
  0.003745,   0.003745,    0.003745,    0.003745,
  0.003683,   0.003683,    0.003683,    0.003683,
  0.003696,   0.003696,    0.003696,    0.003696,
  0.00376,    0.00376,     0.00376,     0.00376,
  0.003794,   0.003794,    0.003794,    0.003794,
  0.00382,    0.00382,     0.00382,     0.00382,
  0.003913,   0.003913,    0.003913,    0.003913,
  0.00393,    0.00393,     0.00393,     0.00393,
  0.003753,   0.003753,    0.003753,    0.003753,
  0.003558,   0.003558,    0.003558,    0.003558,
  0.003501,   0.003501,    0.003501,    0.003501,
  0.003513,   0.003513,    0.003513,    0.003513,
  0.003682,   0.003682,    0.003682,    0.003682,
  0.003899,   0.003899,    0.003899,    0.003899,
  0.003757,   0.003757,    0.003757,    0.003757,
  0.003455,   0.003455,    0.003455,    0.003455,
  0.003404,   0.003404,    0.003404,    0.003404,
  0.00375,    0.00375,     0.00375,     0.00375,
  0.004214,   0.004214,    0.004214,    0.004214,
  0.004354,   0.004354,    0.004354,    0.004354,
  0.004343,   0.004343,    0.004343,    0.004343,
  0.00426,    0.00426,     0.00426,     0.00426,
  0.004185,   0.004185,    0.004185,    0.004185,
  0.00407,    0.00407,     0.00407,     0.00407,
  0.003941,   0.003941,    0.003941,    0.003941,
  0.00384,    0.00384,     0.00384,     0.00384,
  0.00365,    0.00365,     0.00365,     0.00365,
  0.003631,   0.003631,    0.003631,    0.003631,
  0.003645,   0.003645,    0.003645,    0.003645,
  0.00357,    0.00357,     0.00357,     0.00357,
  0.00355,    0.00355,     0.00355,     0.00355,
  0.003812,   0.003812,    0.003812,    0.003812,
  0.004165,   0.004165,    0.004165,    0.004165,
  0.004298,   0.004298,    0.004298,    0.004298,
  0.004305,   0.004305,    0.004305,    0.004305,
  0.004319,   0.004319,    0.004319,    0.004319,
  0.00435,    0.00435,     0.00435,     0.00435,
  0.004367,   0.004367,    0.004367,    0.004367,
  0.004354,   0.004354,    0.004354,    0.004354,
  0.00436,    0.00436,     0.00436,     0.00436,
  0.004385,   0.004385,    0.004385,    0.004385,
  0.004393,   0.004393,    0.004393,    0.004393,
  0.004385,   0.004385,    0.004385,    0.004385,
  0.00436,    0.00436,     0.00436,     0.00436,
  0.004378,   0.004378,    0.004378,    0.004378,
  0.004368,   0.004368,    0.004368,    0.004368,
  0.004318,   0.004318,    0.004318,    0.004318,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004309,   0.004309,    0.004309,    0.004309,
  0.004442,   0.004442,    0.004442,    0.004442,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004511,   0.004511,    0.004511,    0.004511,
  0.004437,   0.004437,    0.004437,    0.004437,
  0.004382,   0.004382,    0.004382,    0.004382,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004196,   0.004196,    0.004196,    0.004196,
  0.004087,   0.004087,    0.004087,    0.004087,
  0.003972,   0.003972,    0.003972,    0.003972,
  0.003861,   0.003861,    0.003861,    0.003861,
  0.003849,   0.003849,    0.003849,    0.003849,
  0.004048,   0.004048,    0.004048,    0.004048,
  0.004249,   0.004249,    0.004249,    0.004249,
  0.00459,    0.00459,     0.00459,     0.00459,
  0.005146,   0.005146,    0.005146,    0.005146,
  0.005349,   0.005349,    0.005349,    0.005349,
  0.005271,   0.005271,    0.005271,    0.005271,
  0.00527,    0.00527,     0.00527,     0.00527,
  0.00516,    0.00516,     0.00516,     0.00516,
  0.005054,   0.005054,    0.005054,    0.005054,
  0.004953,   0.004953,    0.004953,    0.004953,
  0.004959,   0.004959,    0.004959,    0.004959,
  0.005369,   0.005369,    0.005369,    0.005369,
  0.005685,   0.005685,    0.005685,    0.005685,
  0.005695,   0.005695,    0.005695,    0.005695,
  0.005617,   0.005617,    0.005617,    0.005617,
  0.005609,   0.005609,    0.005609,    0.005609,
  0.005761,   0.005761,    0.005761,    0.005761,
  0.005839,   0.005839,    0.005839,    0.005839,
  0.005785,   0.005785,    0.005785,    0.005785,
  0.005762,   0.005762,    0.005762,    0.005762,
  0.005767,   0.005767,    0.005767,    0.005767,
  0.005767,   0.005767,    0.005767,    0.005767,
  0.005789,   0.005789,    0.005789,    0.005789,
  0.005825,   0.005825,    0.005825,    0.005825,
  0.005771,   0.005771,    0.005771,    0.005771,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005435,   0.005435,    0.005435,    0.005435,
  0.005285,   0.005285,    0.005285,    0.005285,
  0.005155,   0.005155,    0.005155,    0.005155,
  0.005051,   0.005051,    0.005051,    0.005051,
  0.005033,   0.005033,    0.005033,    0.005033,
  0.005109,   0.005109,    0.005109,    0.005109,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005536,   0.005536,    0.005536,    0.005536,
  0.005582,   0.005582,    0.005582,    0.005582,
  0.005631,   0.005631,    0.005631,    0.005631,
  0.0057,     0.0057,      0.0057,      0.0057,
  0.005787,   0.005787,    0.005787,    0.005787,
  0.005907,   0.005907,    0.005907,    0.005907,
  0.005996,   0.005996,    0.005996,    0.005996,
  0.006111,   0.006111,    0.006111,    0.006111,
  0.006279,   0.006279,    0.006279,    0.006279,
  0.006293,   0.006293,    0.006293,    0.006293,
  0.005986,   0.005986,    0.005986,    0.005986,
  0.00594,    0.00594,     0.00594,     0.00594,
  0.006134,   0.006134,    0.006134,    0.006134,
  0.005967,   0.005967,    0.005967,    0.005967,
  0.006014,   0.006014,    0.006014,    0.006014,
  0.006231,   0.006231,    0.006231,    0.006231,
  0.006046,   0.006046,    0.006046,    0.006046,
  0.005948,   0.005948,    0.005948,    0.005948,
  0.005989,   0.005989,    0.005989,    0.005989,
  0.005758,   0.005758,    0.005758,    0.005758,
  0.005468,   0.005468,    0.005468,    0.005468,
  0.005394,   0.005394,    0.005394,    0.005394,
  0.005487,   0.005487,    0.005487,    0.005487,
  0.005567,   0.005567,    0.005567,    0.005567,
  0.005486,   0.005486,    0.005486,    0.005486,
  0.005286,   0.005286,    0.005286,    0.005286,
  0.005208,   0.005208,    0.005208,    0.005208,
  0.005288,   0.005288,    0.005288,    0.005288,
  0.005024,   0.005024,    0.005024,    0.005024,
  0.004636,   0.004636,    0.004636,    0.004636,
  0.00452,    0.00452,     0.00452,     0.00452,
  0.004563,   0.004563,    0.004563,    0.004563,
  0.004733,   0.004733,    0.004733,    0.004733,
  0.004848,   0.004848,    0.004848,    0.004848,
  0.004898,   0.004898,    0.004898,    0.004898,
  0.004926,   0.004926,    0.004926,    0.004926,
  0.00502,    0.00502,     0.00502,     0.00502,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005433,   0.005433,    0.005433,    0.005433,
  0.005546,   0.005546,    0.005546,    0.005546,
  0.005622,   0.005622,    0.005622,    0.005622,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005578,   0.005578,    0.005578,    0.005578,
  0.005554,   0.005554,    0.005554,    0.005554,
  0.00547,    0.00547,     0.00547,     0.00547,
  0.005456,   0.005456,    0.005456,    0.005456,
  0.005501,   0.005501,    0.005501,    0.005501,
  0.00555,    0.00555,     0.00555,     0.00555,
  0.005582,   0.005582,    0.005582,    0.005582,
  0.005636,   0.005636,    0.005636,    0.005636,
  0.005732,   0.005732,    0.005732,    0.005732,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.00583,    0.00583,     0.00583,     0.00583,
  0.005874,   0.005874,    0.005874,    0.005874,
  0.005894,   0.005894,    0.005894,    0.005894,
  0.005912,   0.005912,    0.005912,    0.005912,
  0.005931,   0.005931,    0.005931,    0.005931,
  0.005874,   0.005874,    0.005874,    0.005874,
  0.005743,   0.005743,    0.005743,    0.005743,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005438,   0.005438,    0.005438,    0.005438,
  0.005376,   0.005376,    0.005376,    0.005376,
  0.005843,   0.005843,    0.005843,    0.005843,
  0.00618,    0.00618,     0.00618,     0.00618,
  0.005857,   0.005857,    0.005857,    0.005857,
  0.005518,   0.005518,    0.005518,    0.005518,
  0.005279,   0.005279,    0.005279,    0.005279,
  0.005068,   0.005068,    0.005068,    0.005068,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004875,   0.004875,    0.004875,    0.004875,
  0.004906,   0.004906,    0.004906,    0.004906,
  0.004901,   0.004901,    0.004901,    0.004901,
  0.004973,   0.004973,    0.004973,    0.004973,
  0.005049,   0.005049,    0.005049,    0.005049,
  0.005031,   0.005031,    0.005031,    0.005031,
  0.005139,   0.005139,    0.005139,    0.005139,
  0.005355,   0.005355,    0.005355,    0.005355,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005663,   0.005663,    0.005663,    0.005663,
  0.005724,   0.005724,    0.005724,    0.005724,
  0.005778,   0.005778,    0.005778,    0.005778,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.006376,   0.006376,    0.006376,    0.006376,
  0.007053,   0.007053,    0.007053,    0.007053,
  0.007312,   0.007312,    0.007312,    0.007312,
  0.007217,   0.007217,    0.007217,    0.007217,
  0.007232,   0.007232,    0.007232,    0.007232,
  0.007411,   0.007411,    0.007411,    0.007411,
  0.007465,   0.007465,    0.007465,    0.007465,
  0.007386,   0.007386,    0.007386,    0.007386,
  0.00732,    0.00732,     0.00732,     0.00732,
  0.007329,   0.007329,    0.007329,    0.007329,
  0.007349,   0.007349,    0.007349,    0.007349,
  0.007368,   0.007368,    0.007368,    0.007368,
  0.007356,   0.007356,    0.007356,    0.007356,
  0.007313,   0.007313,    0.007313,    0.007313,
  0.007292,   0.007292,    0.007292,    0.007292,
  0.007282,   0.007282,    0.007282,    0.007282,
  0.007272,   0.007272,    0.007272,    0.007272,
  0.007315,   0.007315,    0.007315,    0.007315,
  0.007383,   0.007383,    0.007383,    0.007383,
  0.007408,   0.007408,    0.007408,    0.007408,
  0.007329,   0.007329,    0.007329,    0.007329,
  0.007218,   0.007218,    0.007218,    0.007218,
  0.007089,   0.007089,    0.007089,    0.007089,
  0.006883,   0.006883,    0.006883,    0.006883,
  0.006725,   0.006725,    0.006725,    0.006725,
  0.006681,   0.006681,    0.006681,    0.006681,
  0.006657,   0.006657,    0.006657,    0.006657,
  0.00668,    0.00668,     0.00668,     0.00668,
  0.006712,   0.006712,    0.006712,    0.006712,
  0.006738,   0.006738,    0.006738,    0.006738,
  0.006671,   0.006671,    0.006671,    0.006671,
  0.006386,   0.006386,    0.006386,    0.006386,
  0.006435,   0.006435,    0.006435,    0.006435,
  0.00666,    0.00666,     0.00666,     0.00666,
  0.00675,    0.00675,     0.00675,     0.00675,
  0.006876,   0.006876,    0.006876,    0.006876,
  0.007168,   0.007168,    0.007168,    0.007168,
  0.007453,   0.007453,    0.007453,    0.007453,
  0.007273,   0.007273,    0.007273,    0.007273,
  0.006872,   0.006872,    0.006872,    0.006872,
  0.006967,   0.006967,    0.006967,    0.006967,
  0.007454,   0.007454,    0.007454,    0.007454,
  0.007435,   0.007435,    0.007435,    0.007435,
  0.007209,   0.007209,    0.007209,    0.007209,
  0.00723,    0.00723,     0.00723,     0.00723,
  0.007274,   0.007274,    0.007274,    0.007274,
  0.007339,   0.007339,    0.007339,    0.007339,
  0.007431,   0.007431,    0.007431,    0.007431,
  0.007501,   0.007501,    0.007501,    0.007501,
  0.007515,   0.007515,    0.007515,    0.007515,
  0.007498,   0.007498,    0.007498,    0.007498,
  0.007403,   0.007403,    0.007403,    0.007403,
  0.007286,   0.007286,    0.007286,    0.007286,
  0.007259,   0.007259,    0.007259,    0.007259,
  0.007295,   0.007295,    0.007295,    0.007295,
  0.007272,   0.007272,    0.007272,    0.007272,
  0.007121,   0.007121,    0.007121,    0.007121,
  0.006959,   0.006959,    0.006959,    0.006959,
  0.006851,   0.006851,    0.006851,    0.006851,
  0.006736,   0.006736,    0.006736,    0.006736,
  0.006601,   0.006601,    0.006601,    0.006601,
  0.006518,   0.006518,    0.006518,    0.006518,
  0.00654,    0.00654,     0.00654,     0.00654,
  0.006572,   0.006572,    0.006572,    0.006572,
  0.006507,   0.006507,    0.006507,    0.006507,
  0.00641,    0.00641,     0.00641,     0.00641,
  0.006325,   0.006325,    0.006325,    0.006325,
  0.006298,   0.006298,    0.006298,    0.006298,
  0.006297,   0.006297,    0.006297,    0.006297,
  0.006238,   0.006238,    0.006238,    0.006238,
  0.006195,   0.006195,    0.006195,    0.006195,
  0.006172,   0.006172,    0.006172,    0.006172,
  0.006103,   0.006103,    0.006103,    0.006103,
  0.006055,   0.006055,    0.006055,    0.006055,
  0.005925,   0.005925,    0.005925,    0.005925,
  0.005761,   0.005761,    0.005761,    0.005761,
  0.005657,   0.005657,    0.005657,    0.005657,
  0.005511,   0.005511,    0.005511,    0.005511,
  0.005379,   0.005379,    0.005379,    0.005379,
  0.00515,    0.00515,     0.00515,     0.00515,
  0.004829,   0.004829,    0.004829,    0.004829,
  0.00464,    0.00464,     0.00464,     0.00464,
  0.004507,   0.004507,    0.004507,    0.004507,
  0.004377,   0.004377,    0.004377,    0.004377,
  0.004237,   0.004237,    0.004237,    0.004237,
  0.004143,   0.004143,    0.004143,    0.004143,
  0.003972,   0.003972,    0.003972,    0.003972,
  0.003729,   0.003729,    0.003729,    0.003729,
  0.003577,   0.003577,    0.003577,    0.003577,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.005403,   0.005403,    0.005403,    0.005403,
  0.005917,   0.005917,    0.005917,    0.005917,
  0.005901,   0.005901,    0.005901,    0.005901,
  0.005912,   0.005912,    0.005912,    0.005912,
  0.005896,   0.005896,    0.005896,    0.005896,
  0.005862,   0.005862,    0.005862,    0.005862,
  0.005825,   0.005825,    0.005825,    0.005825,
  0.005804,   0.005804,    0.005804,    0.005804,
  0.005811,   0.005811,    0.005811,    0.005811,
  0.005814,   0.005814,    0.005814,    0.005814,
  0.005811,   0.005811,    0.005811,    0.005811,
  0.005811,   0.005811,    0.005811,    0.005811,
  0.005806,   0.005806,    0.005806,    0.005806,
  0.005806,   0.005806,    0.005806,    0.005806,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.005764,   0.005764,    0.005764,    0.005764,
  0.00573,    0.00573,     0.00573,     0.00573,
  0.005739,   0.005739,    0.005739,    0.005739,
  0.005753,   0.005753,    0.005753,    0.005753,
  0.005771,   0.005771,    0.005771,    0.005771,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.005775,   0.005775,    0.005775,    0.005775,
  0.00583,    0.00583,     0.00583,     0.00583,
  0.005932,   0.005932,    0.005932,    0.005932,
  0.006005,   0.006005,    0.006005,    0.006005,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.005926,   0.005926,    0.005926,    0.005926,
  0.005569,   0.005569,    0.005569,    0.005569,
  0.005291,   0.005291,    0.005291,    0.005291,
  0.005282,   0.005282,    0.005282,    0.005282,
  0.005244,   0.005244,    0.005244,    0.005244,
  0.004946,   0.004946,    0.004946,    0.004946,
  0.004663,   0.004663,    0.004663,    0.004663,
  0.004429,   0.004429,    0.004429,    0.004429,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.00452,    0.00452,     0.00452,     0.00452,
  0.004513,   0.004513,    0.004513,    0.004513,
  0.003986,   0.003986,    0.003986,    0.003986,
  0.003487,   0.003487,    0.003487,    0.003487,
  0.003434,   0.003434,    0.003434,    0.003434,
  0.003475,   0.003475,    0.003475,    0.003475,
  0.003418,   0.003418,    0.003418,    0.003418,
  0.003431,   0.003431,    0.003431,    0.003431,
  0.003614,   0.003614,    0.003614,    0.003614,
  0.003851,   0.003851,    0.003851,    0.003851,
  0.00404,    0.00404,     0.00404,     0.00404,
  0.004413,   0.004413,    0.004413,    0.004413,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004744,   0.004744,    0.004744,    0.004744,
  0.004989,   0.004989,    0.004989,    0.004989,
  0.005239,   0.005239,    0.005239,    0.005239,
  0.005402,   0.005402,    0.005402,    0.005402,
  0.005672,   0.005672,    0.005672,    0.005672,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006211,   0.006211,    0.006211,    0.006211,
  0.006292,   0.006292,    0.006292,    0.006292,
  0.006424,   0.006424,    0.006424,    0.006424,
  0.006536,   0.006536,    0.006536,    0.006536,
  0.006633,   0.006633,    0.006633,    0.006633,
  0.00662,    0.00662,     0.00662,     0.00662,
  0.006563,   0.006563,    0.006563,    0.006563,
  0.006547,   0.006547,    0.006547,    0.006547,
  0.006515,   0.006515,    0.006515,    0.006515,
  0.006508,   0.006508,    0.006508,    0.006508,
  0.006563,   0.006563,    0.006563,    0.006563,
  0.006619,   0.006619,    0.006619,    0.006619,
  0.00664,    0.00664,     0.00664,     0.00664,
  0.006739,   0.006739,    0.006739,    0.006739,
  0.007044,   0.007044,    0.007044,    0.007044,
  0.007266,   0.007266,    0.007266,    0.007266,
  0.007305,   0.007305,    0.007305,    0.007305,
  0.007368,   0.007368,    0.007368,    0.007368,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.007642,   0.007642,    0.007642,    0.007642,
  0.007776,   0.007776,    0.007776,    0.007776,
  0.007821,   0.007821,    0.007821,    0.007821,
  0.007844,   0.007844,    0.007844,    0.007844,
  0.007867,   0.007867,    0.007867,    0.007867,
  0.007813,   0.007813,    0.007813,    0.007813,
  0.007673,   0.007673,    0.007673,    0.007673,
  0.007587,   0.007587,    0.007587,    0.007587,
  0.007551,   0.007551,    0.007551,    0.007551,
  0.007524,   0.007524,    0.007524,    0.007524,
  0.007565,   0.007565,    0.007565,    0.007565,
  0.007444,   0.007444,    0.007444,    0.007444,
  0.007271,   0.007271,    0.007271,    0.007271,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.00725,    0.00725,     0.00725,     0.00725,
  0.007378,   0.007378,    0.007378,    0.007378,
  0.007465,   0.007465,    0.007465,    0.007465,
  0.007499,   0.007499,    0.007499,    0.007499,
  0.007471,   0.007471,    0.007471,    0.007471,
  0.007386,   0.007386,    0.007386,    0.007386,
  0.007274,   0.007274,    0.007274,    0.007274,
  0.007229,   0.007229,    0.007229,    0.007229,
  0.007229,   0.007229,    0.007229,    0.007229,
  0.007208,   0.007208,    0.007208,    0.007208,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007133,   0.007133,    0.007133,    0.007133,
  0.007019,   0.007019,    0.007019,    0.007019,
  0.006717,   0.006717,    0.006717,    0.006717,
  0.006116,   0.006116,    0.006116,    0.006116,
  0.005646,   0.005646,    0.005646,    0.005646,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005412,   0.005412,    0.005412,    0.005412,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005141,   0.005141,    0.005141,    0.005141,
  0.005141,   0.005141,    0.005141,    0.005141,
  0.005066,   0.005066,    0.005066,    0.005066,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004968,   0.004968,    0.004968,    0.004968,
  0.005187,   0.005187,    0.005187,    0.005187,
  0.005743,   0.005743,    0.005743,    0.005743,
  0.006428,   0.006428,    0.006428,    0.006428,
  0.006656,   0.006656,    0.006656,    0.006656,
  0.006519,   0.006519,    0.006519,    0.006519,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.006677,   0.006677,    0.006677,    0.006677,
  0.006896,   0.006896,    0.006896,    0.006896,
  0.006871,   0.006871,    0.006871,    0.006871,
  0.006694,   0.006694,    0.006694,    0.006694,
  0.006558,   0.006558,    0.006558,    0.006558,
  0.006539,   0.006539,    0.006539,    0.006539,
  0.00656,    0.00656,     0.00656,     0.00656,
  0.006596,   0.006596,    0.006596,    0.006596,
  0.006663,   0.006663,    0.006663,    0.006663,
  0.00667,    0.00667,     0.00667,     0.00667,
  0.006643,   0.006643,    0.006643,    0.006643,
  0.006695,   0.006695,    0.006695,    0.006695,
  0.006779,   0.006779,    0.006779,    0.006779,
  0.006665,   0.006665,    0.006665,    0.006665,
  0.006373,   0.006373,    0.006373,    0.006373,
  0.006246,   0.006246,    0.006246,    0.006246,
  0.006277,   0.006277,    0.006277,    0.006277,
  0.006278,   0.006278,    0.006278,    0.006278,
  0.006344,   0.006344,    0.006344,    0.006344,
  0.006573,   0.006573,    0.006573,    0.006573,
  0.006876,   0.006876,    0.006876,    0.006876,
  0.007127,   0.007127,    0.007127,    0.007127,
  0.007236,   0.007236,    0.007236,    0.007236,
  0.007318,   0.007318,    0.007318,    0.007318,
  0.007457,   0.007457,    0.007457,    0.007457,
  0.007502,   0.007502,    0.007502,    0.007502,
  0.007506,   0.007506,    0.007506,    0.007506,
  0.007556,   0.007556,    0.007556,    0.007556,
  0.007607,   0.007607,    0.007607,    0.007607,
  0.007634,   0.007634,    0.007634,    0.007634,
  0.007687,   0.007687,    0.007687,    0.007687,
  0.007739,   0.007739,    0.007739,    0.007739,
  0.007769,   0.007769,    0.007769,    0.007769,
  0.007808,   0.007808,    0.007808,    0.007808,
  0.007856,   0.007856,    0.007856,    0.007856,
  0.007856,   0.007856,    0.007856,    0.007856,
  0.007863,   0.007863,    0.007863,    0.007863,
  0.007895,   0.007895,    0.007895,    0.007895,
  0.007919,   0.007919,    0.007919,    0.007919,
  0.007943,   0.007943,    0.007943,    0.007943,
  0.007991,   0.007991,    0.007991,    0.007991,
  0.008058,   0.008058,    0.008058,    0.008058,
  0.008118,   0.008118,    0.008118,    0.008118,
  0.008188,   0.008188,    0.008188,    0.008188,
  0.008258,   0.008258,    0.008258,    0.008258,
  0.00831,    0.00831,     0.00831,     0.00831,
  0.008386,   0.008386,    0.008386,    0.008386,
  0.008475,   0.008475,    0.008475,    0.008475,
  0.008488,   0.008488,    0.008488,    0.008488,
  0.008528,   0.008528,    0.008528,    0.008528,
  0.008587,   0.008587,    0.008587,    0.008587,
  0.00857,    0.00857,     0.00857,     0.00857,
  0.008608,   0.008608,    0.008608,    0.008608,
  0.008825,   0.008825,    0.008825,    0.008825,
  0.009025,   0.009025,    0.009025,    0.009025,
  0.009106,   0.009106,    0.009106,    0.009106,
  0.009174,   0.009174,    0.009174,    0.009174,
  0.009286,   0.009286,    0.009286,    0.009286,
  0.009371,   0.009371,    0.009371,    0.009371,
  0.009406,   0.009406,    0.009406,    0.009406,
  0.009411,   0.009411,    0.009411,    0.009411,
  0.009433,   0.009433,    0.009433,    0.009433,
  0.009455,   0.009455,    0.009455,    0.009455,
  0.009446,   0.009446,    0.009446,    0.009446,
  0.009466,   0.009466,    0.009466,    0.009466,
  0.009537,   0.009537,    0.009537,    0.009537,
  0.009653,   0.009653,    0.009653,    0.009653,
  0.009818,   0.009818,    0.009818,    0.009818,
  0.00999,    0.00999,     0.00999,     0.00999,
  0.01007,    0.01007,     0.01007,     0.01007,
  0.01017,    0.01017,     0.01017,     0.01017,
  0.01035,    0.01035,     0.01035,     0.01035,
  0.01054,    0.01054,     0.01054,     0.01054,
  0.01068,    0.01068,     0.01068,     0.01068,
  0.01068,    0.01068,     0.01068,     0.01068,
  0.01067,    0.01067,     0.01067,     0.01067,
  0.0106,     0.0106,      0.0106,      0.0106,
  0.01051,    0.01051,     0.01051,     0.01051,
  0.01053,    0.01053,     0.01053,     0.01053,
  0.0105,     0.0105,      0.0105,      0.0105,
  0.01041,    0.01041,     0.01041,     0.01041,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.01008,    0.01008,     0.01008,     0.01008,
  0.009761,   0.009761,    0.009761,    0.009761,
  0.009712,   0.009712,    0.009712,    0.009712,
  0.009838,   0.009838,    0.009838,    0.009838,
  0.009764,   0.009764,    0.009764,    0.009764,
  0.009739,   0.009739,    0.009739,    0.009739,
  0.009843,   0.009843,    0.009843,    0.009843,
  0.01012,    0.01012,     0.01012,     0.01012,
  0.01029,    0.01029,     0.01029,     0.01029,
  0.009968,   0.009968,    0.009968,    0.009968,
  0.009438,   0.009438,    0.009438,    0.009438,
  0.009079,   0.009079,    0.009079,    0.009079,
  0.008676,   0.008676,    0.008676,    0.008676,
  0.00825,    0.00825,     0.00825,     0.00825,
  0.008291,   0.008291,    0.008291,    0.008291,
  0.008265,   0.008265,    0.008265,    0.008265,
  0.008197,   0.008197,    0.008197,    0.008197,
  0.007882,   0.007882,    0.007882,    0.007882,
  0.007204,   0.007204,    0.007204,    0.007204,
  0.006756,   0.006756,    0.006756,    0.006756,
  0.006546,   0.006546,    0.006546,    0.006546,
  0.006308,   0.006308,    0.006308,    0.006308,
  0.005592,   0.005592,    0.005592,    0.005592,
  0.005245,   0.005245,    0.005245,    0.005245,
  0.005405,   0.005405,    0.005405,    0.005405,
  0.005264,   0.005264,    0.005264,    0.005264,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.0039,     0.0039,      0.0039,      0.0039,
  0.003809,   0.003809,    0.003809,    0.003809,
  0.003777,   0.003777,    0.003777,    0.003777,
  0.003872,   0.003872,    0.003872,    0.003872,
  0.004078,   0.004078,    0.004078,    0.004078,
  0.005136,   0.005136,    0.005136,    0.005136,
  0.006886,   0.006886,    0.006886,    0.006886,
  0.007753,   0.007753,    0.007753,    0.007753,
  0.007721,   0.007721,    0.007721,    0.007721,
  0.007807,   0.007807,    0.007807,    0.007807,
  0.008646,   0.008646,    0.008646,    0.008646,
  0.009099,   0.009099,    0.009099,    0.009099,
  0.008419,   0.008419,    0.008419,    0.008419,
  0.00802,    0.00802,     0.00802,     0.00802,
  0.008023,   0.008023,    0.008023,    0.008023,
  0.008032,   0.008032,    0.008032,    0.008032,
  0.008456,   0.008456,    0.008456,    0.008456,
  0.00868,    0.00868,     0.00868,     0.00868,
  0.008507,   0.008507,    0.008507,    0.008507,
  0.008562,   0.008562,    0.008562,    0.008562,
  0.008677,   0.008677,    0.008677,    0.008677,
  0.00874,    0.00874,     0.00874,     0.00874,
  0.00886,    0.00886,     0.00886,     0.00886,
  0.008929,   0.008929,    0.008929,    0.008929,
  0.009007,   0.009007,    0.009007,    0.009007,
  0.008992,   0.008992,    0.008992,    0.008992,
  0.008999,   0.008999,    0.008999,    0.008999,
  0.009065,   0.009065,    0.009065,    0.009065,
  0.009119,   0.009119,    0.009119,    0.009119,
  0.009131,   0.009131,    0.009131,    0.009131,
  0.009023,   0.009023,    0.009023,    0.009023,
  0.008892,   0.008892,    0.008892,    0.008892,
  0.008834,   0.008834,    0.008834,    0.008834,
  0.008879,   0.008879,    0.008879,    0.008879,
  0.008911,   0.008911,    0.008911,    0.008911,
  0.009016,   0.009016,    0.009016,    0.009016,
  0.009126,   0.009126,    0.009126,    0.009126,
  0.009038,   0.009038,    0.009038,    0.009038,
  0.009179,   0.009179,    0.009179,    0.009179,
  0.009205,   0.009205,    0.009205,    0.009205,
  0.009025,   0.009025,    0.009025,    0.009025,
  0.009104,   0.009104,    0.009104,    0.009104,
  0.009028,   0.009028,    0.009028,    0.009028,
  0.008956,   0.008956,    0.008956,    0.008956,
  0.009227,   0.009227,    0.009227,    0.009227,
  0.00961,    0.00961,     0.00961,     0.00961,
  0.00987,    0.00987,     0.00987,     0.00987,
  0.009855,   0.009855,    0.009855,    0.009855,
  0.00978,    0.00978,     0.00978,     0.00978,
  0.009769,   0.009769,    0.009769,    0.009769,
  0.00976,    0.00976,     0.00976,     0.00976,
  0.009631,   0.009631,    0.009631,    0.009631,
  0.009631,   0.009631,    0.009631,    0.009631,
  0.009728,   0.009728,    0.009728,    0.009728,
  0.009639,   0.009639,    0.009639,    0.009639,
  0.009576,   0.009576,    0.009576,    0.009576,
  0.009614,   0.009614,    0.009614,    0.009614,
  0.009759,   0.009759,    0.009759,    0.009759,
  0.00982,    0.00982,     0.00982,     0.00982,
  0.009664,   0.009664,    0.009664,    0.009664,
  0.009558,   0.009558,    0.009558,    0.009558,
  0.009562,   0.009562,    0.009562,    0.009562,
  0.009508,   0.009508,    0.009508,    0.009508,
  0.009401,   0.009401,    0.009401,    0.009401,
  0.009321,   0.009321,    0.009321,    0.009321,
  0.009321,   0.009321,    0.009321,    0.009321,
  0.009401,   0.009401,    0.009401,    0.009401,
  0.009536,   0.009536,    0.009536,    0.009536,
  0.009644,   0.009644,    0.009644,    0.009644,
  0.009617,   0.009617,    0.009617,    0.009617,
  0.009508,   0.009508,    0.009508,    0.009508,
  0.009428,   0.009428,    0.009428,    0.009428,
  0.009321,   0.009321,    0.009321,    0.009321,
  0.009189,   0.009189,    0.009189,    0.009189,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.009059,   0.009059,    0.009059,    0.009059,
  0.009111,   0.009111,    0.009111,    0.009111,
  0.009163,   0.009163,    0.009163,    0.009163,
  0.009322,   0.009322,    0.009322,    0.009322,
  0.009414,   0.009414,    0.009414,    0.009414,
  0.009385,   0.009385,    0.009385,    0.009385,
  0.009337,   0.009337,    0.009337,    0.009337,
  0.009257,   0.009257,    0.009257,    0.009257,
  0.009064,   0.009064,    0.009064,    0.009064,
  0.008721,   0.008721,    0.008721,    0.008721,
  0.008485,   0.008485,    0.008485,    0.008485,
  0.008293,   0.008293,    0.008293,    0.008293,
  0.007922,   0.007922,    0.007922,    0.007922,
  0.007584,   0.007584,    0.007584,    0.007584,
  0.007436,   0.007436,    0.007436,    0.007436,
  0.007363,   0.007363,    0.007363,    0.007363,
  0.007178,   0.007178,    0.007178,    0.007178,
  0.006882,   0.006882,    0.006882,    0.006882,
  0.006694,   0.006694,    0.006694,    0.006694,
  0.0065,     0.0065,      0.0065,      0.0065,
  0.005925,   0.005925,    0.005925,    0.005925,
  0.005435,   0.005435,    0.005435,    0.005435,
  0.005391,   0.005391,    0.005391,    0.005391,
  0.005271,   0.005271,    0.005271,    0.005271,
  0.005146,   0.005146,    0.005146,    0.005146,
  0.005204,   0.005204,    0.005204,    0.005204,
  0.005403,   0.005403,    0.005403,    0.005403,
  0.005617,   0.005617,    0.005617,    0.005617,
  0.006159,   0.006159,    0.006159,    0.006159,
  0.007341,   0.007341,    0.007341,    0.007341,
  0.008559,   0.008559,    0.008559,    0.008559,
  0.009113,   0.009113,    0.009113,    0.009113,
  0.009137,   0.009137,    0.009137,    0.009137,
  0.009095,   0.009095,    0.009095,    0.009095,
  0.009043,   0.009043,    0.009043,    0.009043,
  0.009043,   0.009043,    0.009043,    0.009043,
  0.009106,   0.009106,    0.009106,    0.009106,
  0.009137,   0.009137,    0.009137,    0.009137,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.008855,   0.008855,    0.008855,    0.008855,
  0.008829,   0.008829,    0.008829,    0.008829,
  0.008931,   0.008931,    0.008931,    0.008931,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.008931,   0.008931,    0.008931,    0.008931,
  0.008829,   0.008829,    0.008829,    0.008829,
  0.008778,   0.008778,    0.008778,    0.008778,
  0.008753,   0.008753,    0.008753,    0.008753,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008804,   0.008804,    0.008804,    0.008804,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.009137,   0.009137,    0.009137,    0.009137,
  0.00916,    0.00916,     0.00916,     0.00916,
  0.00913,    0.00913,     0.00913,     0.00913,
  0.009035,   0.009035,    0.009035,    0.009035,
  0.008934,   0.008934,    0.008934,    0.008934,
  0.008759,   0.008759,    0.008759,    0.008759,
  0.00852,    0.00852,     0.00852,     0.00852,
  0.008476,   0.008476,    0.008476,    0.008476,
  0.008398,   0.008398,    0.008398,    0.008398,
  0.007699,   0.007699,    0.007699,    0.007699,
  0.006989,   0.006989,    0.006989,    0.006989,
  0.006972,   0.006972,    0.006972,    0.006972,
  0.006781,   0.006781,    0.006781,    0.006781,
  0.006793,   0.006793,    0.006793,    0.006793,
  0.007498,   0.007498,    0.007498,    0.007498,
  0.00798,    0.00798,     0.00798,     0.00798,
  0.008116,   0.008116,    0.008116,    0.008116,
  0.008224,   0.008224,    0.008224,    0.008224,
  0.008355,   0.008355,    0.008355,    0.008355,
  0.008424,   0.008424,    0.008424,    0.008424,
  0.008358,   0.008358,    0.008358,    0.008358,
  0.008232,   0.008232,    0.008232,    0.008232,
  0.008183,   0.008183,    0.008183,    0.008183,
  0.00834,    0.00834,     0.00834,     0.00834,
  0.008572,   0.008572,    0.008572,    0.008572,
  0.008573,   0.008573,    0.008573,    0.008573,
  0.008079,   0.008079,    0.008079,    0.008079,
  0.007641,   0.007641,    0.007641,    0.007641,
  0.007538,   0.007538,    0.007538,    0.007538,
  0.007373,   0.007373,    0.007373,    0.007373,
  0.007242,   0.007242,    0.007242,    0.007242,
  0.007155,   0.007155,    0.007155,    0.007155,
  0.007133,   0.007133,    0.007133,    0.007133,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007401,   0.007401,    0.007401,    0.007401,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007575,   0.007575,    0.007575,    0.007575,
  0.007465,   0.007465,    0.007465,    0.007465,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007753,   0.007753,    0.007753,    0.007753,
  0.007708,   0.007708,    0.007708,    0.007708,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007708,   0.007708,    0.007708,    0.007708,
  0.007776,   0.007776,    0.007776,    0.007776,
  0.007799,   0.007799,    0.007799,    0.007799,
  0.007776,   0.007776,    0.007776,    0.007776,
  0.007821,   0.007821,    0.007821,    0.007821,
  0.00789,    0.00789,     0.00789,     0.00789,
  0.007951,   0.007951,    0.007951,    0.007951,
  0.007909,   0.007909,    0.007909,    0.007909,
  0.007887,   0.007887,    0.007887,    0.007887,
  0.007946,   0.007946,    0.007946,    0.007946,
  0.007919,   0.007919,    0.007919,    0.007919,
  0.00765,    0.00765,     0.00765,     0.00765,
  0.007313,   0.007313,    0.007313,    0.007313,
  0.007323,   0.007323,    0.007323,    0.007323,
  0.007798,   0.007798,    0.007798,    0.007798,
  0.008044,   0.008044,    0.008044,    0.008044,
  0.00802,    0.00802,     0.00802,     0.00802,
  0.0081,     0.0081,      0.0081,      0.0081,
  0.007997,   0.007997,    0.007997,    0.007997,
  0.007936,   0.007936,    0.007936,    0.007936,
  0.00781,    0.00781,     0.00781,     0.00781,
  0.007516,   0.007516,    0.007516,    0.007516,
  0.007282,   0.007282,    0.007282,    0.007282,
  0.007085,   0.007085,    0.007085,    0.007085,
  0.006788,   0.006788,    0.006788,    0.006788,
  0.006505,   0.006505,    0.006505,    0.006505,
  0.00634,    0.00634,     0.00634,     0.00634,
  0.006248,   0.006248,    0.006248,    0.006248,
  0.006239,   0.006239,    0.006239,    0.006239,
  0.006274,   0.006274,    0.006274,    0.006274,
  0.006277,   0.006277,    0.006277,    0.006277,
  0.006281,   0.006281,    0.006281,    0.006281,
  0.006349,   0.006349,    0.006349,    0.006349,
  0.006455,   0.006455,    0.006455,    0.006455,
  0.006538,   0.006538,    0.006538,    0.006538,
  0.006577,   0.006577,    0.006577,    0.006577,
  0.006616,   0.006616,    0.006616,    0.006616,
  0.006655,   0.006655,    0.006655,    0.006655,
  0.006695,   0.006695,    0.006695,    0.006695,
  0.006715,   0.006715,    0.006715,    0.006715,
  0.006715,   0.006715,    0.006715,    0.006715,
  0.006715,   0.006715,    0.006715,    0.006715,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006775,   0.006775,    0.006775,    0.006775,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006978,   0.006978,    0.006978,    0.006978,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007313,   0.007313,    0.007313,    0.007313,
  0.0074,     0.0074,      0.0074,      0.0074,
  0.007418,   0.007418,    0.007418,    0.007418,
  0.007304,   0.007304,    0.007304,    0.007304,
  0.007291,   0.007291,    0.007291,    0.007291,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007017,   0.007017,    0.007017,    0.007017,
  0.006901,   0.006901,    0.006901,    0.006901,
  0.006787,   0.006787,    0.006787,    0.006787,
  0.006624,   0.006624,    0.006624,    0.006624,
  0.006534,   0.006534,    0.006534,    0.006534,
  0.006493,   0.006493,    0.006493,    0.006493,
  0.006394,   0.006394,    0.006394,    0.006394,
  0.006368,   0.006368,    0.006368,    0.006368,
  0.006301,   0.006301,    0.006301,    0.006301,
  0.006175,   0.006175,    0.006175,    0.006175,
  0.006152,   0.006152,    0.006152,    0.006152,
  0.006161,   0.006161,    0.006161,    0.006161,
  0.006161,   0.006161,    0.006161,    0.006161,
  0.006203,   0.006203,    0.006203,    0.006203,
  0.006341,   0.006341,    0.006341,    0.006341,
  0.006435,   0.006435,    0.006435,    0.006435,
  0.006444,   0.006444,    0.006444,    0.006444,
  0.006472,   0.006472,    0.006472,    0.006472,
  0.006451,   0.006451,    0.006451,    0.006451,
  0.006337,   0.006337,    0.006337,    0.006337,
  0.006268,   0.006268,    0.006268,    0.006268,
  0.006286,   0.006286,    0.006286,    0.006286,
  0.006313,   0.006313,    0.006313,    0.006313,
  0.006204,   0.006204,    0.006204,    0.006204,
  0.006026,   0.006026,    0.006026,    0.006026,
  0.005893,   0.005893,    0.005893,    0.005893,
  0.005837,   0.005837,    0.005837,    0.005837,
  0.0058,     0.0058,      0.0058,      0.0058,
  0.005719,   0.005719,    0.005719,    0.005719,
  0.005682,   0.005682,    0.005682,    0.005682,
  0.005654,   0.005654,    0.005654,    0.005654,
  0.005582,   0.005582,    0.005582,    0.005582,
  0.005542,   0.005542,    0.005542,    0.005542,
  0.005497,   0.005497,    0.005497,    0.005497,
  0.005439,   0.005439,    0.005439,    0.005439,
  0.005422,   0.005422,    0.005422,    0.005422,
  0.00537,    0.00537,     0.00537,     0.00537,
  0.005351,   0.005351,    0.005351,    0.005351,
  0.005489,   0.005489,    0.005489,    0.005489,
  0.005608,   0.005608,    0.005608,    0.005608,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005175,   0.005175,    0.005175,    0.005175,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004456,   0.004456,    0.004456,    0.004456,
  0.00454,    0.00454,     0.00454,     0.00454,
  0.004803,   0.004803,    0.004803,    0.004803,
  0.004805,   0.004805,    0.004805,    0.004805,
  0.004589,   0.004589,    0.004589,    0.004589,
  0.004599,   0.004599,    0.004599,    0.004599,
  0.004616,   0.004616,    0.004616,    0.004616,
  0.004531,   0.004531,    0.004531,    0.004531,
  0.004182,   0.004182,    0.004182,    0.004182,
  0.003784,   0.003784,    0.003784,    0.003784,
  0.004036,   0.004036,    0.004036,    0.004036,
  0.00413,    0.00413,     0.00413,     0.00413,
  0.004153,   0.004153,    0.004153,    0.004153,
  0.004319,   0.004319,    0.004319,    0.004319,
  0.004256,   0.004256,    0.004256,    0.004256,
  0.004209,   0.004209,    0.004209,    0.004209,
  0.004145,   0.004145,    0.004145,    0.004145,
  0.004161,   0.004161,    0.004161,    0.004161,
  0.004107,   0.004107,    0.004107,    0.004107,
  0.003984,   0.003984,    0.003984,    0.003984,
  0.003992,   0.003992,    0.003992,    0.003992,
  0.003981,   0.003981,    0.003981,    0.003981,
  0.003986,   0.003986,    0.003986,    0.003986,
  0.00405,    0.00405,     0.00405,     0.00405,
  0.004256,   0.004256,    0.004256,    0.004256,
  0.004572,   0.004572,    0.004572,    0.004572,
  0.004741,   0.004741,    0.004741,    0.004741,
  0.004737,   0.004737,    0.004737,    0.004737,
  0.004723,   0.004723,    0.004723,    0.004723,
  0.004728,   0.004728,    0.004728,    0.004728,
  0.004733,   0.004733,    0.004733,    0.004733,
  0.00473,    0.00473,     0.00473,     0.00473,
  0.00465,    0.00465,     0.00465,     0.00465,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004477,   0.004477,    0.004477,    0.004477,
  0.004398,   0.004398,    0.004398,    0.004398,
  0.004384,   0.004384,    0.004384,    0.004384,
  0.004358,   0.004358,    0.004358,    0.004358,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004418,   0.004418,    0.004418,    0.004418,
  0.004434,   0.004434,    0.004434,    0.004434,
  0.004495,   0.004495,    0.004495,    0.004495,
  0.004604,   0.004604,    0.004604,    0.004604,
  0.004702,   0.004702,    0.004702,    0.004702,
  0.004669,   0.004669,    0.004669,    0.004669,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004368,   0.004368,    0.004368,    0.004368,
  0.004153,   0.004153,    0.004153,    0.004153,
  0.003911,   0.003911,    0.003911,    0.003911,
  0.003728,   0.003728,    0.003728,    0.003728,
  0.00364,    0.00364,     0.00364,     0.00364,
  0.003628,   0.003628,    0.003628,    0.003628,
  0.003648,   0.003648,    0.003648,    0.003648,
  0.003629,   0.003629,    0.003629,    0.003629,
  0.003578,   0.003578,    0.003578,    0.003578,
  0.003531,   0.003531,    0.003531,    0.003531,
  0.003439,   0.003439,    0.003439,    0.003439,
  0.003368,   0.003368,    0.003368,    0.003368,
  0.00331,    0.00331,     0.00331,     0.00331,
  0.003202,   0.003202,    0.003202,    0.003202,
  0.003088,   0.003088,    0.003088,    0.003088,
  0.003017,   0.003017,    0.003017,    0.003017,
  0.003035,   0.003035,    0.003035,    0.003035,
  0.003097,   0.003097,    0.003097,    0.003097,
  0.003134,   0.003134,    0.003134,    0.003134,
  0.00319,    0.00319,     0.00319,     0.00319,
  0.003374,   0.003374,    0.003374,    0.003374,
  0.003475,   0.003475,    0.003475,    0.003475,
  0.003664,   0.003664,    0.003664,    0.003664,
  0.00397,    0.00397,     0.00397,     0.00397,
  0.004146,   0.004146,    0.004146,    0.004146,
  0.004429,   0.004429,    0.004429,    0.004429,
  0.004655,   0.004655,    0.004655,    0.004655,
  0.004718,   0.004718,    0.004718,    0.004718,
  0.004806,   0.004806,    0.004806,    0.004806,
  0.004981,   0.004981,    0.004981,    0.004981,
  0.005125,   0.005125,    0.005125,    0.005125,
  0.005191,   0.005191,    0.005191,    0.005191,
  0.005204,   0.005204,    0.005204,    0.005204,
  0.005192,   0.005192,    0.005192,    0.005192,
  0.005187,   0.005187,    0.005187,    0.005187,
  0.005186,   0.005186,    0.005186,    0.005186,
  0.005195,   0.005195,    0.005195,    0.005195,
  0.005196,   0.005196,    0.005196,    0.005196,
  0.005167,   0.005167,    0.005167,    0.005167,
  0.005161,   0.005161,    0.005161,    0.005161,
  0.005158,   0.005158,    0.005158,    0.005158,
  0.00509,    0.00509,     0.00509,     0.00509,
  0.005021,   0.005021,    0.005021,    0.005021,
  0.004971,   0.004971,    0.004971,    0.004971,
  0.004949,   0.004949,    0.004949,    0.004949,
  0.005014,   0.005014,    0.005014,    0.005014,
  0.005093,   0.005093,    0.005093,    0.005093,
  0.005043,   0.005043,    0.005043,    0.005043,
  0.004621,   0.004621,    0.004621,    0.004621,
  0.004099,   0.004099,    0.004099,    0.004099,
  0.003681,   0.003681,    0.003681,    0.003681,
  0.003298,   0.003298,    0.003298,    0.003298,
  0.003084,   0.003084,    0.003084,    0.003084,
  0.002946,   0.002946,    0.002946,    0.002946,
  0.002889,   0.002889,    0.002889,    0.002889,
  0.002934,   0.002934,    0.002934,    0.002934,
  0.002958,   0.002958,    0.002958,    0.002958,
  0.002891,   0.002891,    0.002891,    0.002891,
  0.002835,   0.002835,    0.002835,    0.002835,
  0.002845,   0.002845,    0.002845,    0.002845,
  0.002726,   0.002726,    0.002726,    0.002726,
  0.002446,   0.002446,    0.002446,    0.002446,
  0.002358,   0.002358,    0.002358,    0.002358,
  0.00229,    0.00229,     0.00229,     0.00229,
  0.002224,   0.002224,    0.002224,    0.002224,
  0.002402,   0.002402,    0.002402,    0.002402,
  0.002495,   0.002495,    0.002495,    0.002495,
  0.002443,   0.002443,    0.002443,    0.002443,
  0.002447,   0.002447,    0.002447,    0.002447,
  0.002711,   0.002711,    0.002711,    0.002711,
  0.003037,   0.003037,    0.003037,    0.003037,
  0.00376,    0.00376,     0.00376,     0.00376,
  0.004964,   0.004964,    0.004964,    0.004964,
  0.005562,   0.005562,    0.005562,    0.005562,
  0.005612,   0.005612,    0.005612,    0.005612,
  0.005615,   0.005615,    0.005615,    0.005615,
  0.005538,   0.005538,    0.005538,    0.005538,
  0.005476,   0.005476,    0.005476,    0.005476,
  0.00548,    0.00548,     0.00548,     0.00548,
  0.005471,   0.005471,    0.005471,    0.005471,
  0.005383,   0.005383,    0.005383,    0.005383,
  0.005308,   0.005308,    0.005308,    0.005308,
  0.00525,    0.00525,     0.00525,     0.00525,
  0.00519,    0.00519,     0.00519,     0.00519,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005207,   0.005207,    0.005207,    0.005207,
  0.005219,   0.005219,    0.005219,    0.005219,
  0.005155,   0.005155,    0.005155,    0.005155,
  0.005123,   0.005123,    0.005123,    0.005123,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.004996,   0.004996,    0.004996,    0.004996,
  0.005076,   0.005076,    0.005076,    0.005076,
  0.005061,   0.005061,    0.005061,    0.005061,
  0.005076,   0.005076,    0.005076,    0.005076,
  0.005394,   0.005394,    0.005394,    0.005394,
  0.005605,   0.005605,    0.005605,    0.005605,
  0.005618,   0.005618,    0.005618,    0.005618,
  0.005578,   0.005578,    0.005578,    0.005578,
  0.005244,   0.005244,    0.005244,    0.005244,
  0.004789,   0.004789,    0.004789,    0.004789,
  0.004622,   0.004622,    0.004622,    0.004622,
  0.004686,   0.004686,    0.004686,    0.004686,
  0.00454,    0.00454,     0.00454,     0.00454,
  0.004177,   0.004177,    0.004177,    0.004177,
  0.004234,   0.004234,    0.004234,    0.004234,
  0.004585,   0.004585,    0.004585,    0.004585,
  0.004693,   0.004693,    0.004693,    0.004693,
  0.004665,   0.004665,    0.004665,    0.004665,
  0.004725,   0.004725,    0.004725,    0.004725,
  0.004644,   0.004644,    0.004644,    0.004644,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.004002,   0.004002,    0.004002,    0.004002,
  0.004118,   0.004118,    0.004118,    0.004118,
  0.003961,   0.003961,    0.003961,    0.003961,
  0.003908,   0.003908,    0.003908,    0.003908,
  0.00371,    0.00371,     0.00371,     0.00371,
  0.003389,   0.003389,    0.003389,    0.003389,
  0.003407,   0.003407,    0.003407,    0.003407,
  0.003457,   0.003457,    0.003457,    0.003457,
  0.003488,   0.003488,    0.003488,    0.003488,
  0.003633,   0.003633,    0.003633,    0.003633,
  0.004042,   0.004042,    0.004042,    0.004042,
  0.004677,   0.004677,    0.004677,    0.004677,
  0.005146,   0.005146,    0.005146,    0.005146,
  0.005468,   0.005468,    0.005468,    0.005468,
  0.005918,   0.005918,    0.005918,    0.005918,
  0.006409,   0.006409,    0.006409,    0.006409,
  0.00684,    0.00684,     0.00684,     0.00684,
  0.007169,   0.007169,    0.007169,    0.007169,
  0.007209,   0.007209,    0.007209,    0.007209,
  0.007156,   0.007156,    0.007156,    0.007156,
  0.007182,   0.007182,    0.007182,    0.007182,
  0.007135,   0.007135,    0.007135,    0.007135,
  0.007039,   0.007039,    0.007039,    0.007039,
  0.006924,   0.006924,    0.006924,    0.006924,
  0.006767,   0.006767,    0.006767,    0.006767,
  0.00662,    0.00662,     0.00662,     0.00662,
  0.006474,   0.006474,    0.006474,    0.006474,
  0.006348,   0.006348,    0.006348,    0.006348,
  0.006242,   0.006242,    0.006242,    0.006242,
  0.00617,    0.00617,     0.00617,     0.00617,
  0.006108,   0.006108,    0.006108,    0.006108,
  0.006197,   0.006197,    0.006197,    0.006197,
  0.006251,   0.006251,    0.006251,    0.006251,
  0.006122,   0.006122,    0.006122,    0.006122,
  0.005994,   0.005994,    0.005994,    0.005994,
  0.005855,   0.005855,    0.005855,    0.005855,
  0.005811,   0.005811,    0.005811,    0.005811,
  0.005664,   0.005664,    0.005664,    0.005664,
  0.005423,   0.005423,    0.005423,    0.005423,
  0.005371,   0.005371,    0.005371,    0.005371,
  0.005445,   0.005445,    0.005445,    0.005445,
  0.005437,   0.005437,    0.005437,    0.005437,
  0.005439,   0.005439,    0.005439,    0.005439,
  0.005578,   0.005578,    0.005578,    0.005578,
  0.005723,   0.005723,    0.005723,    0.005723,
  0.005764,   0.005764,    0.005764,    0.005764,
  0.005694,   0.005694,    0.005694,    0.005694,
  0.005663,   0.005663,    0.005663,    0.005663,
  0.005638,   0.005638,    0.005638,    0.005638,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.005096,   0.005096,    0.005096,    0.005096,
  0.004964,   0.004964,    0.004964,    0.004964,
  0.004982,   0.004982,    0.004982,    0.004982,
  0.004894,   0.004894,    0.004894,    0.004894,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004868,   0.004868,    0.004868,    0.004868,
  0.004919,   0.004919,    0.004919,    0.004919,
  0.005065,   0.005065,    0.005065,    0.005065,
  0.004898,   0.004898,    0.004898,    0.004898,
  0.004732,   0.004732,    0.004732,    0.004732,
  0.004819,   0.004819,    0.004819,    0.004819,
  0.004936,   0.004936,    0.004936,    0.004936,
  0.004865,   0.004865,    0.004865,    0.004865,
  0.004836,   0.004836,    0.004836,    0.004836,
  0.004872,   0.004872,    0.004872,    0.004872,
  0.004718,   0.004718,    0.004718,    0.004718,
  0.004517,   0.004517,    0.004517,    0.004517,
  0.004411,   0.004411,    0.004411,    0.004411,
  0.004403,   0.004403,    0.004403,    0.004403,
  0.004553,   0.004553,    0.004553,    0.004553,
  0.00481,    0.00481,     0.00481,     0.00481,
  0.004942,   0.004942,    0.004942,    0.004942,
  0.004891,   0.004891,    0.004891,    0.004891,
  0.004784,   0.004784,    0.004784,    0.004784,
  0.004765,   0.004765,    0.004765,    0.004765,
  0.00481,    0.00481,     0.00481,     0.00481,
  0.004798,   0.004798,    0.004798,    0.004798,
  0.004803,   0.004803,    0.004803,    0.004803,
  0.004904,   0.004904,    0.004904,    0.004904,
  0.005026,   0.005026,    0.005026,    0.005026,
  0.005124,   0.005124,    0.005124,    0.005124,
  0.005203,   0.005203,    0.005203,    0.005203,
  0.005259,   0.005259,    0.005259,    0.005259,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005355,   0.005355,    0.005355,    0.005355,
  0.005423,   0.005423,    0.005423,    0.005423,
  0.005455,   0.005455,    0.005455,    0.005455,
  0.005464,   0.005464,    0.005464,    0.005464,
  0.005487,   0.005487,    0.005487,    0.005487,
  0.005374,   0.005374,    0.005374,    0.005374,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005101,   0.005101,    0.005101,    0.005101,
  0.005058,   0.005058,    0.005058,    0.005058,
  0.005069,   0.005069,    0.005069,    0.005069,
  0.005062,   0.005062,    0.005062,    0.005062,
  0.0051,     0.0051,      0.0051,      0.0051,
  0.005244,   0.005244,    0.005244,    0.005244,
  0.00537,    0.00537,     0.00537,     0.00537,
  0.005389,   0.005389,    0.005389,    0.005389,
  0.005377,   0.005377,    0.005377,    0.005377,
  0.005334,   0.005334,    0.005334,    0.005334,
  0.005379,   0.005379,    0.005379,    0.005379,
  0.005437,   0.005437,    0.005437,    0.005437,
  0.005435,   0.005435,    0.005435,    0.005435,
  0.005579,   0.005579,    0.005579,    0.005579,
  0.005702,   0.005702,    0.005702,    0.005702,
  0.005779,   0.005779,    0.005779,    0.005779,
  0.005876,   0.005876,    0.005876,    0.005876,
  0.005949,   0.005949,    0.005949,    0.005949,
  0.005952,   0.005952,    0.005952,    0.005952,
  0.005912,   0.005912,    0.005912,    0.005912,
  0.005837,   0.005837,    0.005837,    0.005837,
  0.005743,   0.005743,    0.005743,    0.005743,
  0.005672,   0.005672,    0.005672,    0.005672,
  0.005641,   0.005641,    0.005641,    0.005641,
  0.005615,   0.005615,    0.005615,    0.005615,
  0.005542,   0.005542,    0.005542,    0.005542,
  0.005471,   0.005471,    0.005471,    0.005471,
  0.005433,   0.005433,    0.005433,    0.005433,
  0.005364,   0.005364,    0.005364,    0.005364,
  0.005282,   0.005282,    0.005282,    0.005282,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005107,   0.005107,    0.005107,    0.005107,
  0.005155,   0.005155,    0.005155,    0.005155,
  0.005346,   0.005346,    0.005346,    0.005346,
  0.005511,   0.005511,    0.005511,    0.005511,
  0.005808,   0.005808,    0.005808,    0.005808,
  0.00601,    0.00601,     0.00601,     0.00601,
  0.005881,   0.005881,    0.005881,    0.005881,
  0.00567,    0.00567,     0.00567,     0.00567,
  0.005592,   0.005592,    0.005592,    0.005592,
  0.005601,   0.005601,    0.005601,    0.005601,
  0.005593,   0.005593,    0.005593,    0.005593,
  0.005528,   0.005528,    0.005528,    0.005528,
  0.00549,    0.00549,     0.00549,     0.00549,
  0.005454,   0.005454,    0.005454,    0.005454,
  0.005468,   0.005468,    0.005468,    0.005468,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005405,   0.005405,    0.005405,    0.005405,
  0.005376,   0.005376,    0.005376,    0.005376,
  0.005061,   0.005061,    0.005061,    0.005061,
  0.004601,   0.004601,    0.004601,    0.004601,
  0.004286,   0.004286,    0.004286,    0.004286,
  0.004122,   0.004122,    0.004122,    0.004122,
  0.004066,   0.004066,    0.004066,    0.004066,
  0.004146,   0.004146,    0.004146,    0.004146,
  0.004317,   0.004317,    0.004317,    0.004317,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.00447,    0.00447,     0.00447,     0.00447,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.003494,   0.003494,    0.003494,    0.003494,
  0.0033,     0.0033,      0.0033,      0.0033,
  0.004025,   0.004025,    0.004025,    0.004025,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.005142,   0.005142,    0.005142,    0.005142,
  0.005469,   0.005469,    0.005469,    0.005469,
  0.005678,   0.005678,    0.005678,    0.005678,
  0.005874,   0.005874,    0.005874,    0.005874,
  0.006054,   0.006054,    0.006054,    0.006054,
  0.006194,   0.006194,    0.006194,    0.006194,
  0.006262,   0.006262,    0.006262,    0.006262,
  0.006282,   0.006282,    0.006282,    0.006282,
  0.006272,   0.006272,    0.006272,    0.006272,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006283,   0.006283,    0.006283,    0.006283,
  0.006321,   0.006321,    0.006321,    0.006321,
  0.006359,   0.006359,    0.006359,    0.006359,
  0.006359,   0.006359,    0.006359,    0.006359,
  0.006359,   0.006359,    0.006359,    0.006359,
  0.006391,   0.006391,    0.006391,    0.006391,
  0.006334,   0.006334,    0.006334,    0.006334,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006177,   0.006177,    0.006177,    0.006177,
  0.006022,   0.006022,    0.006022,    0.006022,
  0.005911,   0.005911,    0.005911,    0.005911,
  0.005773,   0.005773,    0.005773,    0.005773,
  0.005696,   0.005696,    0.005696,    0.005696,
  0.005708,   0.005708,    0.005708,    0.005708,
  0.005743,   0.005743,    0.005743,    0.005743,
  0.005779,   0.005779,    0.005779,    0.005779,
  0.00578,    0.00578,     0.00578,     0.00578,
  0.005633,   0.005633,    0.005633,    0.005633,
  0.005337,   0.005337,    0.005337,    0.005337,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.004791,   0.004791,    0.004791,    0.004791,
  0.004409,   0.004409,    0.004409,    0.004409,
  0.004033,   0.004033,    0.004033,    0.004033,
  0.003513,   0.003513,    0.003513,    0.003513,
  0.003131,   0.003131,    0.003131,    0.003131,
  0.003064,   0.003064,    0.003064,    0.003064,
  0.003003,   0.003003,    0.003003,    0.003003,
  0.003006,   0.003006,    0.003006,    0.003006,
  0.00301,    0.00301,     0.00301,     0.00301,
  0.002984,   0.002984,    0.002984,    0.002984,
  0.003017,   0.003017,    0.003017,    0.003017,
  0.003108,   0.003108,    0.003108,    0.003108,
  0.003296,   0.003296,    0.003296,    0.003296,
  0.003419,   0.003419,    0.003419,    0.003419,
  0.003478,   0.003478,    0.003478,    0.003478,
  0.003538,   0.003538,    0.003538,    0.003538,
  0.0036,     0.0036,      0.0036,      0.0036,
  0.003641,   0.003641,    0.003641,    0.003641,
  0.003832,   0.003832,    0.003832,    0.003832,
  0.004147,   0.004147,    0.004147,    0.004147,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004556,   0.004556,    0.004556,    0.004556,
  0.004658,   0.004658,    0.004658,    0.004658,
  0.004704,   0.004704,    0.004704,    0.004704,
  0.004819,   0.004819,    0.004819,    0.004819,
  0.004883,   0.004883,    0.004883,    0.004883,
  0.004924,   0.004924,    0.004924,    0.004924,
  0.004919,   0.004919,    0.004919,    0.004919,
  0.004845,   0.004845,    0.004845,    0.004845,
  0.004751,   0.004751,    0.004751,    0.004751,
  0.004628,   0.004628,    0.004628,    0.004628,
  0.004475,   0.004475,    0.004475,    0.004475,
  0.004313,   0.004313,    0.004313,    0.004313,
  0.004195,   0.004195,    0.004195,    0.004195,
  0.00413,    0.00413,     0.00413,     0.00413,
  0.00411,    0.00411,     0.00411,     0.00411,
  0.004105,   0.004105,    0.004105,    0.004105,
  0.004048,   0.004048,    0.004048,    0.004048,
  0.004005,   0.004005,    0.004005,    0.004005,
  0.004051,   0.004051,    0.004051,    0.004051,
  0.003757,   0.003757,    0.003757,    0.003757,
  0.003192,   0.003192,    0.003192,    0.003192,
  0.00274,    0.00274,     0.00274,     0.00274,
  0.002448,   0.002448,    0.002448,    0.002448,
  0.002423,   0.002423,    0.002423,    0.002423,
  0.002493,   0.002493,    0.002493,    0.002493,
  0.002341,   0.002341,    0.002341,    0.002341,
  0.002155,   0.002155,    0.002155,    0.002155,
  0.002228,   0.002228,    0.002228,    0.002228,
  0.002244,   0.002244,    0.002244,    0.002244,
  0.002201,   0.002201,    0.002201,    0.002201,
  0.002283,   0.002283,    0.002283,    0.002283,
  0.002406,   0.002406,    0.002406,    0.002406,
  0.00256,    0.00256,     0.00256,     0.00256,
  0.002616,   0.002616,    0.002616,    0.002616,
  0.002614,   0.002614,    0.002614,    0.002614,
  0.002609,   0.002609,    0.002609,    0.002609,
  0.002605,   0.002605,    0.002605,    0.002605,
  0.002666,   0.002666,    0.002666,    0.002666,
  0.002668,   0.002668,    0.002668,    0.002668,
  0.002611,   0.002611,    0.002611,    0.002611,
  0.002656,   0.002656,    0.002656,    0.002656,
  0.002731,   0.002731,    0.002731,    0.002731,
  0.002773,   0.002773,    0.002773,    0.002773,
  0.002852,   0.002852,    0.002852,    0.002852,
  0.002956,   0.002956,    0.002956,    0.002956,
  0.003166,   0.003166,    0.003166,    0.003166,
  0.003432,   0.003432,    0.003432,    0.003432,
  0.003636,   0.003636,    0.003636,    0.003636,
  0.003886,   0.003886,    0.003886,    0.003886,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.00451,    0.00451,     0.00451,     0.00451,
  0.004591,   0.004591,    0.004591,    0.004591,
  0.004503,   0.004503,    0.004503,    0.004503,
  0.004331,   0.004331,    0.004331,    0.004331,
  0.004104,   0.004104,    0.004104,    0.004104,
  0.0039,     0.0039,      0.0039,      0.0039,
  0.003837,   0.003837,    0.003837,    0.003837,
  0.003865,   0.003865,    0.003865,    0.003865,
  0.003947,   0.003947,    0.003947,    0.003947,
  0.004039,   0.004039,    0.004039,    0.004039,
  0.00416,    0.00416,     0.00416,     0.00416,
  0.004246,   0.004246,    0.004246,    0.004246,
  0.004275,   0.004275,    0.004275,    0.004275,
  0.004331,   0.004331,    0.004331,    0.004331,
  0.00431,    0.00431,     0.00431,     0.00431,
  0.004137,   0.004137,    0.004137,    0.004137,
  0.0041,     0.0041,      0.0041,      0.0041,
  0.004203,   0.004203,    0.004203,    0.004203,
  0.004207,   0.004207,    0.004207,    0.004207,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004069,   0.004069,    0.004069,    0.004069,
  0.003982,   0.003982,    0.003982,    0.003982,
  0.003846,   0.003846,    0.003846,    0.003846,
  0.003646,   0.003646,    0.003646,    0.003646,
  0.003472,   0.003472,    0.003472,    0.003472,
  0.003242,   0.003242,    0.003242,    0.003242,
  0.002997,   0.002997,    0.002997,    0.002997,
  0.00289,    0.00289,     0.00289,     0.00289,
  0.002912,   0.002912,    0.002912,    0.002912,
  0.003002,   0.003002,    0.003002,    0.003002,
  0.003098,   0.003098,    0.003098,    0.003098,
  0.003351,   0.003351,    0.003351,    0.003351,
  0.003604,   0.003604,    0.003604,    0.003604,
  0.003702,   0.003702,    0.003702,    0.003702,
  0.003736,   0.003736,    0.003736,    0.003736,
  0.003674,   0.003674,    0.003674,    0.003674,
  0.003611,   0.003611,    0.003611,    0.003611,
  0.003608,   0.003608,    0.003608,    0.003608,
  0.003792,   0.003792,    0.003792,    0.003792,
  0.004072,   0.004072,    0.004072,    0.004072,
  0.004369,   0.004369,    0.004369,    0.004369,
  0.004706,   0.004706,    0.004706,    0.004706,
  0.005007,   0.005007,    0.005007,    0.005007,
  0.005221,   0.005221,    0.005221,    0.005221,
  0.005384,   0.005384,    0.005384,    0.005384,
  0.005346,   0.005346,    0.005346,    0.005346,
  0.004972,   0.004972,    0.004972,    0.004972,
  0.004671,   0.004671,    0.004671,    0.004671,
  0.004738,   0.004738,    0.004738,    0.004738,
  0.004913,   0.004913,    0.004913,    0.004913,
  0.005024,   0.005024,    0.005024,    0.005024,
  0.005157,   0.005157,    0.005157,    0.005157,
  0.005283,   0.005283,    0.005283,    0.005283,
  0.005326,   0.005326,    0.005326,    0.005326,
  0.005319,   0.005319,    0.005319,    0.005319,
  0.005298,   0.005298,    0.005298,    0.005298,
  0.005256,   0.005256,    0.005256,    0.005256,
  0.005172,   0.005172,    0.005172,    0.005172,
  0.005081,   0.005081,    0.005081,    0.005081,
  0.005025,   0.005025,    0.005025,    0.005025,
  0.004953,   0.004953,    0.004953,    0.004953,
  0.004885,   0.004885,    0.004885,    0.004885,
  0.004825,   0.004825,    0.004825,    0.004825,
  0.004793,   0.004793,    0.004793,    0.004793,
  0.004841,   0.004841,    0.004841,    0.004841,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004883,   0.004883,    0.004883,    0.004883,
  0.004882,   0.004882,    0.004882,    0.004882,
  0.004823,   0.004823,    0.004823,    0.004823,
  0.004824,   0.004824,    0.004824,    0.004824,
  0.00484,    0.00484,     0.00484,     0.00484,
  0.004609,   0.004609,    0.004609,    0.004609,
  0.004073,   0.004073,    0.004073,    0.004073,
  0.003541,   0.003541,    0.003541,    0.003541,
  0.00323,    0.00323,     0.00323,     0.00323,
  0.003015,   0.003015,    0.003015,    0.003015,
  0.002896,   0.002896,    0.002896,    0.002896,
  0.002904,   0.002904,    0.002904,    0.002904,
  0.002887,   0.002887,    0.002887,    0.002887,
  0.002898,   0.002898,    0.002898,    0.002898,
  0.00281,    0.00281,     0.00281,     0.00281,
  0.00263,    0.00263,     0.00263,     0.00263,
  0.002539,   0.002539,    0.002539,    0.002539,
  0.002322,   0.002322,    0.002322,    0.002322,
  0.002141,   0.002141,    0.002141,    0.002141,
  0.002169,   0.002169,    0.002169,    0.002169,
  0.002224,   0.002224,    0.002224,    0.002224,
  0.002338,   0.002338,    0.002338,    0.002338,
  0.002471,   0.002471,    0.002471,    0.002471,
  0.00273,    0.00273,     0.00273,     0.00273,
  0.003071,   0.003071,    0.003071,    0.003071,
  0.003314,   0.003314,    0.003314,    0.003314,
  0.003579,   0.003579,    0.003579,    0.003579,
  0.003863,   0.003863,    0.003863,    0.003863,
  0.004118,   0.004118,    0.004118,    0.004118,
  0.004539,   0.004539,    0.004539,    0.004539,
  0.005043,   0.005043,    0.005043,    0.005043,
  0.005302,   0.005302,    0.005302,    0.005302,
  0.005356,   0.005356,    0.005356,    0.005356,
  0.005367,   0.005367,    0.005367,    0.005367,
  0.005366,   0.005366,    0.005366,    0.005366,
  0.00537,    0.00537,     0.00537,     0.00537,
  0.005368,   0.005368,    0.005368,    0.005368,
  0.005317,   0.005317,    0.005317,    0.005317,
  0.00533,    0.00533,     0.00533,     0.00533,
  0.005372,   0.005372,    0.005372,    0.005372,
  0.005358,   0.005358,    0.005358,    0.005358,
  0.005376,   0.005376,    0.005376,    0.005376,
  0.005402,   0.005402,    0.005402,    0.005402,
  0.005357,   0.005357,    0.005357,    0.005357,
  0.005202,   0.005202,    0.005202,    0.005202,
  0.004916,   0.004916,    0.004916,    0.004916,
  0.00463,    0.00463,     0.00463,     0.00463,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.003624,   0.003624,    0.003624,    0.003624,
  0.003229,   0.003229,    0.003229,    0.003229,
  0.003002,   0.003002,    0.003002,    0.003002,
  0.002594,   0.002594,    0.002594,    0.002594,
  0.002222,   0.002222,    0.002222,    0.002222,
  0.00211,    0.00211,     0.00211,     0.00211,
  0.001971,   0.001971,    0.001971,    0.001971,
  0.00189,    0.00189,     0.00189,     0.00189,
  0.00191,    0.00191,     0.00191,     0.00191,
  0.001865,   0.001865,    0.001865,    0.001865,
  0.001765,   0.001765,    0.001765,    0.001765,
  0.001813,   0.001813,    0.001813,    0.001813,
  0.001855,   0.001855,    0.001855,    0.001855,
  0.001838,   0.001838,    0.001838,    0.001838,
  0.001829,   0.001829,    0.001829,    0.001829,
  0.001908,   0.001908,    0.001908,    0.001908,
  0.001934,   0.001934,    0.001934,    0.001934,
  0.001908,   0.001908,    0.001908,    0.001908,
  0.001945,   0.001945,    0.001945,    0.001945,
  0.002023,   0.002023,    0.002023,    0.002023,
  0.002081,   0.002081,    0.002081,    0.002081,
  0.002092,   0.002092,    0.002092,    0.002092,
  0.002264,   0.002264,    0.002264,    0.002264,
  0.002598,   0.002598,    0.002598,    0.002598,
  0.003843,   0.003843,    0.003843,    0.003843,
  0.00533,    0.00533,     0.00533,     0.00533,
  0.005821,   0.005821,    0.005821,    0.005821,
  0.005906,   0.005906,    0.005906,    0.005906,
  0.005967,   0.005967,    0.005967,    0.005967,
  0.005901,   0.005901,    0.005901,    0.005901,
  0.005813,   0.005813,    0.005813,    0.005813,
  0.005818,   0.005818,    0.005818,    0.005818,
  0.005823,   0.005823,    0.005823,    0.005823,
  0.005815,   0.005815,    0.005815,    0.005815,
  0.005854,   0.005854,    0.005854,    0.005854,
  0.005912,   0.005912,    0.005912,    0.005912,
  0.005949,   0.005949,    0.005949,    0.005949,
  0.005981,   0.005981,    0.005981,    0.005981,
  0.005946,   0.005946,    0.005946,    0.005946,
  0.005833,   0.005833,    0.005833,    0.005833,
  0.005745,   0.005745,    0.005745,    0.005745,
  0.005758,   0.005758,    0.005758,    0.005758,
  0.005825,   0.005825,    0.005825,    0.005825,
  0.005983,   0.005983,    0.005983,    0.005983,
  0.006273,   0.006273,    0.006273,    0.006273,
  0.006568,   0.006568,    0.006568,    0.006568,
  0.006718,   0.006718,    0.006718,    0.006718,
  0.006724,   0.006724,    0.006724,    0.006724,
  0.006697,   0.006697,    0.006697,    0.006697,
  0.00649,    0.00649,     0.00649,     0.00649,
  0.006122,   0.006122,    0.006122,    0.006122,
  0.005701,   0.005701,    0.005701,    0.005701,
  0.005198,   0.005198,    0.005198,    0.005198,
  0.005182,   0.005182,    0.005182,    0.005182,
  0.005157,   0.005157,    0.005157,    0.005157,
  0.004979,   0.004979,    0.004979,    0.004979,
  0.005157,   0.005157,    0.005157,    0.005157,
  0.00508,    0.00508,     0.00508,     0.00508,
  0.004732,   0.004732,    0.004732,    0.004732,
  0.004732,   0.004732,    0.004732,    0.004732,
  0.005062,   0.005062,    0.005062,    0.005062,
  0.005068,   0.005068,    0.005068,    0.005068,
  0.004824,   0.004824,    0.004824,    0.004824,
  0.004754,   0.004754,    0.004754,    0.004754,
  0.004654,   0.004654,    0.004654,    0.004654,
  0.004666,   0.004666,    0.004666,    0.004666,
  0.004899,   0.004899,    0.004899,    0.004899,
  0.005208,   0.005208,    0.005208,    0.005208,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005264,   0.005264,    0.005264,    0.005264,
  0.005033,   0.005033,    0.005033,    0.005033,
  0.004938,   0.004938,    0.004938,    0.004938,
  0.005367,   0.005367,    0.005367,    0.005367,
  0.006339,   0.006339,    0.006339,    0.006339,
  0.007168,   0.007168,    0.007168,    0.007168,
  0.00742,    0.00742,     0.00742,     0.00742,
  0.007457,   0.007457,    0.007457,    0.007457,
  0.007589,   0.007589,    0.007589,    0.007589,
  0.007651,   0.007651,    0.007651,    0.007651,
  0.007559,   0.007559,    0.007559,    0.007559,
  0.007437,   0.007437,    0.007437,    0.007437,
  0.007387,   0.007387,    0.007387,    0.007387,
  0.007365,   0.007365,    0.007365,    0.007365,
  0.007347,   0.007347,    0.007347,    0.007347,
  0.007337,   0.007337,    0.007337,    0.007337,
  0.007343,   0.007343,    0.007343,    0.007343,
  0.007342,   0.007342,    0.007342,    0.007342,
  0.007342,   0.007342,    0.007342,    0.007342,
  0.007405,   0.007405,    0.007405,    0.007405,
  0.00746,    0.00746,     0.00746,     0.00746,
  0.007488,   0.007488,    0.007488,    0.007488,
  0.007526,   0.007526,    0.007526,    0.007526,
  0.007559,   0.007559,    0.007559,    0.007559,
  0.007512,   0.007512,    0.007512,    0.007512,
  0.007376,   0.007376,    0.007376,    0.007376,
  0.006837,   0.006837,    0.006837,    0.006837,
  0.005976,   0.005976,    0.005976,    0.005976,
  0.005072,   0.005072,    0.005072,    0.005072,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.003499,   0.003499,    0.003499,    0.003499,
  0.003472,   0.003472,    0.003472,    0.003472,
  0.003341,   0.003341,    0.003341,    0.003341,
  0.002906,   0.002906,    0.002906,    0.002906,
  0.002659,   0.002659,    0.002659,    0.002659,
  0.002486,   0.002486,    0.002486,    0.002486,
  0.002328,   0.002328,    0.002328,    0.002328,
  0.002295,   0.002295,    0.002295,    0.002295,
  0.00234,    0.00234,     0.00234,     0.00234,
  0.002353,   0.002353,    0.002353,    0.002353,
  0.002437,   0.002437,    0.002437,    0.002437,
  0.002531,   0.002531,    0.002531,    0.002531,
  0.002531,   0.002531,    0.002531,    0.002531,
  0.002437,   0.002437,    0.002437,    0.002437,
  0.00229,    0.00229,     0.00229,     0.00229,
  0.002251,   0.002251,    0.002251,    0.002251,
  0.002462,   0.002462,    0.002462,    0.002462,
  0.002714,   0.002714,    0.002714,    0.002714,
  0.002953,   0.002953,    0.002953,    0.002953,
  0.003191,   0.003191,    0.003191,    0.003191,
  0.003351,   0.003351,    0.003351,    0.003351,
  0.003618,   0.003618,    0.003618,    0.003618,
  0.003882,   0.003882,    0.003882,    0.003882,
  0.004055,   0.004055,    0.004055,    0.004055,
  0.004177,   0.004177,    0.004177,    0.004177,
  0.004286,   0.004286,    0.004286,    0.004286,
  0.004465,   0.004465,    0.004465,    0.004465,
  0.004723,   0.004723,    0.004723,    0.004723,
  0.004949,   0.004949,    0.004949,    0.004949,
  0.005151,   0.005151,    0.005151,    0.005151,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005621,   0.005621,    0.005621,    0.005621,
  0.00576,    0.00576,     0.00576,     0.00576,
  0.005806,   0.005806,    0.005806,    0.005806,
  0.005855,   0.005855,    0.005855,    0.005855,
  0.005907,   0.005907,    0.005907,    0.005907,
  0.005896,   0.005896,    0.005896,    0.005896,
  0.005947,   0.005947,    0.005947,    0.005947,
  0.006041,   0.006041,    0.006041,    0.006041,
  0.006036,   0.006036,    0.006036,    0.006036,
  0.005929,   0.005929,    0.005929,    0.005929,
  0.005914,   0.005914,    0.005914,    0.005914,
  0.005969,   0.005969,    0.005969,    0.005969,
  0.005902,   0.005902,    0.005902,    0.005902,
  0.005728,   0.005728,    0.005728,    0.005728,
  0.005617,   0.005617,    0.005617,    0.005617,
  0.00558,    0.00558,     0.00558,     0.00558,
  0.005631,   0.005631,    0.005631,    0.005631,
  0.005676,   0.005676,    0.005676,    0.005676,
  0.005308,   0.005308,    0.005308,    0.005308,
  0.004837,   0.004837,    0.004837,    0.004837,
  0.004638,   0.004638,    0.004638,    0.004638,
  0.004596,   0.004596,    0.004596,    0.004596,
  0.004617,   0.004617,    0.004617,    0.004617,
  0.004249,   0.004249,    0.004249,    0.004249,
  0.00339,    0.00339,     0.00339,     0.00339,
  0.002915,   0.002915,    0.002915,    0.002915,
  0.003055,   0.003055,    0.003055,    0.003055,
  0.003497,   0.003497,    0.003497,    0.003497,
  0.003451,   0.003451,    0.003451,    0.003451,
  0.003325,   0.003325,    0.003325,    0.003325,
  0.003766,   0.003766,    0.003766,    0.003766,
  0.004081,   0.004081,    0.004081,    0.004081,
  0.004272,   0.004272,    0.004272,    0.004272,
  0.004509,   0.004509,    0.004509,    0.004509,
  0.004713,   0.004713,    0.004713,    0.004713,
  0.004841,   0.004841,    0.004841,    0.004841,
  0.005134,   0.005134,    0.005134,    0.005134,
  0.005437,   0.005437,    0.005437,    0.005437,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005986,   0.005986,    0.005986,    0.005986,
  0.006241,   0.006241,    0.006241,    0.006241,
  0.006519,   0.006519,    0.006519,    0.006519,
  0.00668,    0.00668,     0.00668,     0.00668,
  0.006619,   0.006619,    0.006619,    0.006619,
  0.006677,   0.006677,    0.006677,    0.006677,
  0.006863,   0.006863,    0.006863,    0.006863,
  0.007094,   0.007094,    0.007094,    0.007094,
  0.007223,   0.007223,    0.007223,    0.007223,
  0.007308,   0.007308,    0.007308,    0.007308,
  0.007472,   0.007472,    0.007472,    0.007472,
  0.007589,   0.007589,    0.007589,    0.007589,
  0.007551,   0.007551,    0.007551,    0.007551,
  0.007508,   0.007508,    0.007508,    0.007508,
  0.007461,   0.007461,    0.007461,    0.007461,
  0.007387,   0.007387,    0.007387,    0.007387,
  0.00732,    0.00732,     0.00732,     0.00732,
  0.007265,   0.007265,    0.007265,    0.007265,
  0.007178,   0.007178,    0.007178,    0.007178,
  0.007121,   0.007121,    0.007121,    0.007121,
  0.007127,   0.007127,    0.007127,    0.007127,
  0.007146,   0.007146,    0.007146,    0.007146,
  0.007246,   0.007246,    0.007246,    0.007246,
  0.007392,   0.007392,    0.007392,    0.007392,
  0.007425,   0.007425,    0.007425,    0.007425,
  0.007364,   0.007364,    0.007364,    0.007364,
  0.007347,   0.007347,    0.007347,    0.007347,
  0.007271,   0.007271,    0.007271,    0.007271,
  0.007035,   0.007035,    0.007035,    0.007035,
  0.006697,   0.006697,    0.006697,    0.006697,
  0.006489,   0.006489,    0.006489,    0.006489,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006061,   0.006061,    0.006061,    0.006061,
  0.00583,    0.00583,     0.00583,     0.00583,
  0.006114,   0.006114,    0.006114,    0.006114,
  0.006557,   0.006557,    0.006557,    0.006557,
  0.006707,   0.006707,    0.006707,    0.006707,
  0.007684,   0.007684,    0.007684,    0.007684,
  0.009327,   0.009327,    0.009327,    0.009327,
  0.01011,    0.01011,     0.01011,     0.01011,
  0.01048,    0.01048,     0.01048,     0.01048,
  0.01088,    0.01088,     0.01088,     0.01088,
  0.01104,    0.01104,     0.01104,     0.01104,
  0.01104,    0.01104,     0.01104,     0.01104,
  0.01104,    0.01104,     0.01104,     0.01104,
  0.0111,     0.0111,      0.0111,      0.0111,
  0.01119,    0.01119,     0.01119,     0.01119,
  0.01119,    0.01119,     0.01119,     0.01119,
  0.01072,    0.01072,     0.01072,     0.01072,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.01021,    0.01021,     0.01021,     0.01021,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.01016,    0.01016,     0.01016,     0.01016,
  0.01008,    0.01008,     0.01008,     0.01008,
  0.01021,    0.01021,     0.01021,     0.01021,
  0.01028,    0.01028,     0.01028,     0.01028,
  0.01028,    0.01028,     0.01028,     0.01028,
  0.01035,    0.01035,     0.01035,     0.01035,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.0102,     0.0102,      0.0102,      0.0102,
  0.01018,    0.01018,     0.01018,     0.01018,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.01019,    0.01019,     0.01019,     0.01019,
  0.0101,     0.0101,      0.0101,      0.0101,
  0.01007,    0.01007,     0.01007,     0.01007,
  0.01012,    0.01012,     0.01012,     0.01012,
  0.01022,    0.01022,     0.01022,     0.01022,
  0.01028,    0.01028,     0.01028,     0.01028,
  0.01028,    0.01028,     0.01028,     0.01028,
  0.01034,    0.01034,     0.01034,     0.01034,
  0.01046,    0.01046,     0.01046,     0.01046,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.0107,     0.0107,      0.0107,      0.0107,
  0.0107,     0.0107,      0.0107,      0.0107,
  0.01067,    0.01067,     0.01067,     0.01067,
  0.0107,     0.0107,      0.0107,      0.0107,
  0.01082,    0.01082,     0.01082,     0.01082,
  0.01098,    0.01098,     0.01098,     0.01098,
  0.01107,    0.01107,     0.01107,     0.01107,
  0.01088,    0.01088,     0.01088,     0.01088,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01047,    0.01047,     0.01047,     0.01047,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.0107,     0.0107,      0.0107,      0.0107,
  0.01078,    0.01078,     0.01078,     0.01078,
  0.01075,    0.01075,     0.01075,     0.01075,
  0.01072,    0.01072,     0.01072,     0.01072,
  0.009817,   0.009817,    0.009817,    0.009817,
  0.008699,   0.008699,    0.008699,    0.008699,
  0.008198,   0.008198,    0.008198,    0.008198,
  0.007771,   0.007771,    0.007771,    0.007771,
  0.007603,   0.007603,    0.007603,    0.007603,
  0.007539,   0.007539,    0.007539,    0.007539,
  0.007537,   0.007537,    0.007537,    0.007537,
  0.007824,   0.007824,    0.007824,    0.007824,
  0.008344,   0.008344,    0.008344,    0.008344,
  0.008717,   0.008717,    0.008717,    0.008717,
  0.008991,   0.008991,    0.008991,    0.008991,
  0.009039,   0.009039,    0.009039,    0.009039,
  0.008827,   0.008827,    0.008827,    0.008827,
  0.008582,   0.008582,    0.008582,    0.008582,
  0.00839,    0.00839,     0.00839,     0.00839,
  0.008262,   0.008262,    0.008262,    0.008262,
  0.008146,   0.008146,    0.008146,    0.008146,
  0.00809,    0.00809,     0.00809,     0.00809,
  0.00802,    0.00802,     0.00802,     0.00802,
  0.007836,   0.007836,    0.007836,    0.007836,
  0.007708,   0.007708,    0.007708,    0.007708,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007641,   0.007641,    0.007641,    0.007641,
  0.007754,   0.007754,    0.007754,    0.007754,
  0.00796,    0.00796,     0.00796,     0.00796,
  0.008195,   0.008195,    0.008195,    0.008195,
  0.008353,   0.008353,    0.008353,    0.008353,
  0.008451,   0.008451,    0.008451,    0.008451,
  0.008488,   0.008488,    0.008488,    0.008488,
  0.008457,   0.008457,    0.008457,    0.008457,
  0.008408,   0.008408,    0.008408,    0.008408,
  0.00836,    0.00836,     0.00836,     0.00836,
  0.008312,   0.008312,    0.008312,    0.008312,
  0.008267,   0.008267,    0.008267,    0.008267,
  0.008018,   0.008018,    0.008018,    0.008018,
  0.007603,   0.007603,    0.007603,    0.007603,
  0.007444,   0.007444,    0.007444,    0.007444,
  0.007195,   0.007195,    0.007195,    0.007195,
  0.006513,   0.006513,    0.006513,    0.006513,
  0.006088,   0.006088,    0.006088,    0.006088,
  0.00598,    0.00598,     0.00598,     0.00598,
  0.005865,   0.005865,    0.005865,    0.005865,
  0.005694,   0.005694,    0.005694,    0.005694,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005566,   0.005566,    0.005566,    0.005566,
  0.00559,    0.00559,     0.00559,     0.00559,
  0.005637,   0.005637,    0.005637,    0.005637,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005586,   0.005586,    0.005586,    0.005586,
  0.005515,   0.005515,    0.005515,    0.005515,
  0.005385,   0.005385,    0.005385,    0.005385,
  0.005715,   0.005715,    0.005715,    0.005715,
  0.006402,   0.006402,    0.006402,    0.006402,
  0.006816,   0.006816,    0.006816,    0.006816,
  0.006982,   0.006982,    0.006982,    0.006982,
  0.007179,   0.007179,    0.007179,    0.007179,
  0.00733,    0.00733,     0.00733,     0.00733,
  0.007497,   0.007497,    0.007497,    0.007497,
  0.007609,   0.007609,    0.007609,    0.007609,
  0.007475,   0.007475,    0.007475,    0.007475,
  0.007232,   0.007232,    0.007232,    0.007232,
  0.007124,   0.007124,    0.007124,    0.007124,
  0.007178,   0.007178,    0.007178,    0.007178,
  0.007226,   0.007226,    0.007226,    0.007226,
  0.007296,   0.007296,    0.007296,    0.007296,
  0.007413,   0.007413,    0.007413,    0.007413,
  0.0075,     0.0075,      0.0075,      0.0075,
  0.007523,   0.007523,    0.007523,    0.007523,
  0.007516,   0.007516,    0.007516,    0.007516,
  0.007486,   0.007486,    0.007486,    0.007486,
  0.007472,   0.007472,    0.007472,    0.007472,
  0.007503,   0.007503,    0.007503,    0.007503,
  0.007556,   0.007556,    0.007556,    0.007556,
  0.007669,   0.007669,    0.007669,    0.007669,
  0.007782,   0.007782,    0.007782,    0.007782,
  0.007792,   0.007792,    0.007792,    0.007792,
  0.007785,   0.007785,    0.007785,    0.007785,
  0.0078,     0.0078,      0.0078,      0.0078,
  0.007769,   0.007769,    0.007769,    0.007769,
  0.007605,   0.007605,    0.007605,    0.007605,
  0.007367,   0.007367,    0.007367,    0.007367,
  0.007169,   0.007169,    0.007169,    0.007169,
  0.006762,   0.006762,    0.006762,    0.006762,
  0.006359,   0.006359,    0.006359,    0.006359,
  0.006244,   0.006244,    0.006244,    0.006244,
  0.006161,   0.006161,    0.006161,    0.006161,
  0.006148,   0.006148,    0.006148,    0.006148,
  0.006084,   0.006084,    0.006084,    0.006084,
  0.006089,   0.006089,    0.006089,    0.006089,
  0.006168,   0.006168,    0.006168,    0.006168,
  0.006241,   0.006241,    0.006241,    0.006241,
  0.006378,   0.006378,    0.006378,    0.006378,
  0.006352,   0.006352,    0.006352,    0.006352,
  0.006264,   0.006264,    0.006264,    0.006264,
  0.006283,   0.006283,    0.006283,    0.006283,
  0.006262,   0.006262,    0.006262,    0.006262,
  0.006146,   0.006146,    0.006146,    0.006146,
  0.006063,   0.006063,    0.006063,    0.006063,
  0.005974,   0.005974,    0.005974,    0.005974,
  0.006195,   0.006195,    0.006195,    0.006195,
  0.006665,   0.006665,    0.006665,    0.006665,
  0.006932,   0.006932,    0.006932,    0.006932,
  0.006955,   0.006955,    0.006955,    0.006955,
  0.006879,   0.006879,    0.006879,    0.006879,
  0.006958,   0.006958,    0.006958,    0.006958,
  0.007193,   0.007193,    0.007193,    0.007193,
  0.007315,   0.007315,    0.007315,    0.007315,
  0.007296,   0.007296,    0.007296,    0.007296,
  0.007099,   0.007099,    0.007099,    0.007099,
  0.006751,   0.006751,    0.006751,    0.006751,
  0.006624,   0.006624,    0.006624,    0.006624,
  0.006655,   0.006655,    0.006655,    0.006655,
  0.006719,   0.006719,    0.006719,    0.006719,
  0.006848,   0.006848,    0.006848,    0.006848,
  0.006949,   0.006949,    0.006949,    0.006949,
  0.007052,   0.007052,    0.007052,    0.007052,
  0.007152,   0.007152,    0.007152,    0.007152,
  0.007154,   0.007154,    0.007154,    0.007154,
  0.007095,   0.007095,    0.007095,    0.007095,
  0.007095,   0.007095,    0.007095,    0.007095,
  0.007053,   0.007053,    0.007053,    0.007053,
  0.006981,   0.006981,    0.006981,    0.006981,
  0.006942,   0.006942,    0.006942,    0.006942,
  0.00697,    0.00697,     0.00697,     0.00697,
  0.006974,   0.006974,    0.006974,    0.006974,
  0.006887,   0.006887,    0.006887,    0.006887,
  0.006962,   0.006962,    0.006962,    0.006962,
  0.007035,   0.007035,    0.007035,    0.007035,
  0.00705,    0.00705,     0.00705,     0.00705,
  0.007082,   0.007082,    0.007082,    0.007082,
  0.007097,   0.007097,    0.007097,    0.007097,
  0.007116,   0.007116,    0.007116,    0.007116,
  0.007067,   0.007067,    0.007067,    0.007067,
  0.007095,   0.007095,    0.007095,    0.007095,
  0.007398,   0.007398,    0.007398,    0.007398,
  0.00789,    0.00789,     0.00789,     0.00789,
  0.008414,   0.008414,    0.008414,    0.008414,
  0.008507,   0.008507,    0.008507,    0.008507,
  0.008974,   0.008974,    0.008974,    0.008974,
  0.01059,    0.01059,     0.01059,     0.01059,
  0.01174,    0.01174,     0.01174,     0.01174,
  0.01203,    0.01203,     0.01203,     0.01203,
  0.01206,    0.01206,     0.01206,     0.01206,
  0.0119,     0.0119,      0.0119,      0.0119,
  0.0118,     0.0118,      0.0118,      0.0118,
  0.01173,    0.01173,     0.01173,     0.01173,
  0.01167,    0.01167,     0.01167,     0.01167,
  0.01164,    0.01164,     0.01164,     0.01164,
  0.0116,     0.0116,      0.0116,      0.0116,
  0.01154,    0.01154,     0.01154,     0.01154,
  0.01144,    0.01144,     0.01144,     0.01144,
  0.01132,    0.01132,     0.01132,     0.01132,
  0.01125,    0.01125,     0.01125,     0.01125,
  0.01119,    0.01119,     0.01119,     0.01119,
  0.01116,    0.01116,     0.01116,     0.01116,
  0.01119,    0.01119,     0.01119,     0.01119,
  0.01116,    0.01116,     0.01116,     0.01116,
  0.01116,    0.01116,     0.01116,     0.01116,
  0.01113,    0.01113,     0.01113,     0.01113,
  0.01062,    0.01062,     0.01062,     0.01062,
  0.009979,   0.009979,    0.009979,    0.009979,
  0.009645,   0.009645,    0.009645,    0.009645,
  0.009455,   0.009455,    0.009455,    0.009455,
  0.009374,   0.009374,    0.009374,    0.009374,
  0.009348,   0.009348,    0.009348,    0.009348,
  0.009401,   0.009401,    0.009401,    0.009401,
  0.009481,   0.009481,    0.009481,    0.009481,
  0.009481,   0.009481,    0.009481,    0.009481,
  0.009423,   0.009423,    0.009423,    0.009423,
  0.009418,   0.009418,    0.009418,    0.009418,
  0.009382,   0.009382,    0.009382,    0.009382,
  0.009369,   0.009369,    0.009369,    0.009369,
  0.009412,   0.009412,    0.009412,    0.009412,
  0.00944,    0.00944,     0.00944,     0.00944,
  0.009495,   0.009495,    0.009495,    0.009495,
  0.009446,   0.009446,    0.009446,    0.009446,
  0.009346,   0.009346,    0.009346,    0.009346,
  0.009338,   0.009338,    0.009338,    0.009338,
  0.009302,   0.009302,    0.009302,    0.009302,
  0.009218,   0.009218,    0.009218,    0.009218,
  0.009265,   0.009265,    0.009265,    0.009265,
  0.00903,    0.00903,     0.00903,     0.00903,
  0.00849,    0.00849,     0.00849,     0.00849,
  0.008301,   0.008301,    0.008301,    0.008301,
  0.008614,   0.008614,    0.008614,    0.008614,
  0.008975,   0.008975,    0.008975,    0.008975,
  0.008838,   0.008838,    0.008838,    0.008838,
  0.008285,   0.008285,    0.008285,    0.008285,
  0.008177,   0.008177,    0.008177,    0.008177,
  0.008389,   0.008389,    0.008389,    0.008389,
  0.008392,   0.008392,    0.008392,    0.008392,
  0.00836,    0.00836,     0.00836,     0.00836,
  0.008203,   0.008203,    0.008203,    0.008203,
  0.008137,   0.008137,    0.008137,    0.008137,
  0.008133,   0.008133,    0.008133,    0.008133,
  0.007951,   0.007951,    0.007951,    0.007951,
  0.007857,   0.007857,    0.007857,    0.007857,
  0.00806,    0.00806,     0.00806,     0.00806,
  0.008298,   0.008298,    0.008298,    0.008298,
  0.008451,   0.008451,    0.008451,    0.008451,
  0.008515,   0.008515,    0.008515,    0.008515,
  0.00852,    0.00852,     0.00852,     0.00852,
  0.008591,   0.008591,    0.008591,    0.008591,
  0.008633,   0.008633,    0.008633,    0.008633,
  0.00868,    0.00868,     0.00868,     0.00868,
  0.00879,    0.00879,     0.00879,     0.00879,
  0.008896,   0.008896,    0.008896,    0.008896,
  0.008948,   0.008948,    0.008948,    0.008948,
  0.009065,   0.009065,    0.009065,    0.009065,
  0.009212,   0.009212,    0.009212,    0.009212,
  0.009256,   0.009256,    0.009256,    0.009256,
  0.009355,   0.009355,    0.009355,    0.009355,
  0.009401,   0.009401,    0.009401,    0.009401,
  0.009348,   0.009348,    0.009348,    0.009348,
  0.009348,   0.009348,    0.009348,    0.009348,
  0.009321,   0.009321,    0.009321,    0.009321,
  0.009321,   0.009321,    0.009321,    0.009321,
  0.009348,   0.009348,    0.009348,    0.009348,
  0.009401,   0.009401,    0.009401,    0.009401,
  0.009481,   0.009481,    0.009481,    0.009481,
  0.009673,   0.009673,    0.009673,    0.009673,
  0.00981,    0.00981,     0.00981,     0.00981,
  0.009681,   0.009681,    0.009681,    0.009681,
  0.009478,   0.009478,    0.009478,    0.009478,
  0.00915,    0.00915,     0.00915,     0.00915,
  0.008955,   0.008955,    0.008955,    0.008955,
  0.008835,   0.008835,    0.008835,    0.008835,
  0.008593,   0.008593,    0.008593,    0.008593,
  0.008438,   0.008438,    0.008438,    0.008438,
  0.008344,   0.008344,    0.008344,    0.008344,
  0.008394,   0.008394,    0.008394,    0.008394,
  0.008396,   0.008396,    0.008396,    0.008396,
  0.008204,   0.008204,    0.008204,    0.008204,
  0.008127,   0.008127,    0.008127,    0.008127,
  0.008217,   0.008217,    0.008217,    0.008217,
  0.008702,   0.008702,    0.008702,    0.008702,
  0.008866,   0.008866,    0.008866,    0.008866,
  0.009115,   0.009115,    0.009115,    0.009115,
  0.01004,    0.01004,     0.01004,     0.01004,
  0.01045,    0.01045,     0.01045,     0.01045,
  0.01039,    0.01039,     0.01039,     0.01039,
  0.009967,   0.009967,    0.009967,    0.009967,
  0.009587,   0.009587,    0.009587,    0.009587,
  0.009465,   0.009465,    0.009465,    0.009465,
  0.009499,   0.009499,    0.009499,    0.009499,
  0.009689,   0.009689,    0.009689,    0.009689,
  0.009689,   0.009689,    0.009689,    0.009689,
  0.009668,   0.009668,    0.009668,    0.009668,
  0.009748,   0.009748,    0.009748,    0.009748,
  0.009753,   0.009753,    0.009753,    0.009753,
  0.00973,    0.00973,     0.00973,     0.00973,
  0.009694,   0.009694,    0.009694,    0.009694,
  0.009565,   0.009565,    0.009565,    0.009565,
  0.009487,   0.009487,    0.009487,    0.009487,
  0.009468,   0.009468,    0.009468,    0.009468,
  0.00937,    0.00937,     0.00937,     0.00937,
  0.009268,   0.009268,    0.009268,    0.009268,
  0.009216,   0.009216,    0.009216,    0.009216,
  0.009216,   0.009216,    0.009216,    0.009216,
  0.009189,   0.009189,    0.009189,    0.009189,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.008931,   0.008931,    0.008931,    0.008931,
  0.008956,   0.008956,    0.008956,    0.008956,
  0.009008,   0.009008,    0.009008,    0.009008,
  0.009059,   0.009059,    0.009059,    0.009059,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.009122,   0.009122,    0.009122,    0.009122,
  0.00905,    0.00905,     0.00905,     0.00905,
  0.00891,    0.00891,     0.00891,     0.00891,
  0.008838,   0.008838,    0.008838,    0.008838,
  0.008775,   0.008775,    0.008775,    0.008775,
  0.00872,    0.00872,     0.00872,     0.00872,
  0.008797,   0.008797,    0.008797,    0.008797,
  0.008995,   0.008995,    0.008995,    0.008995,
  0.009103,   0.009103,    0.009103,    0.009103,
  0.009087,   0.009087,    0.009087,    0.009087,
  0.008956,   0.008956,    0.008956,    0.008956,
  0.008829,   0.008829,    0.008829,    0.008829,
  0.008956,   0.008956,    0.008956,    0.008956,
  0.009542,   0.009542,    0.009542,    0.009542,
  0.009801,   0.009801,    0.009801,    0.009801,
  0.009511,   0.009511,    0.009511,    0.009511,
  0.0095,     0.0095,      0.0095,      0.0095,
  0.009581,   0.009581,    0.009581,    0.009581,
  0.009597,   0.009597,    0.009597,    0.009597,
  0.009585,   0.009585,    0.009585,    0.009585,
  0.009561,   0.009561,    0.009561,    0.009561,
  0.009428,   0.009428,    0.009428,    0.009428,
  0.009098,   0.009098,    0.009098,    0.009098,
  0.008888,   0.008888,    0.008888,    0.008888,
  0.008665,   0.008665,    0.008665,    0.008665,
  0.008297,   0.008297,    0.008297,    0.008297,
  0.007935,   0.007935,    0.007935,    0.007935,
  0.007634,   0.007634,    0.007634,    0.007634,
  0.007482,   0.007482,    0.007482,    0.007482,
  0.007449,   0.007449,    0.007449,    0.007449,
  0.007415,   0.007415,    0.007415,    0.007415,
  0.007485,   0.007485,    0.007485,    0.007485,
  0.00743,    0.00743,     0.00743,     0.00743,
  0.007311,   0.007311,    0.007311,    0.007311,
  0.007343,   0.007343,    0.007343,    0.007343,
  0.007382,   0.007382,    0.007382,    0.007382,
  0.007452,   0.007452,    0.007452,    0.007452,
  0.007468,   0.007468,    0.007468,    0.007468,
  0.00746,    0.00746,     0.00746,     0.00746,
  0.007476,   0.007476,    0.007476,    0.007476,
  0.007493,   0.007493,    0.007493,    0.007493,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007526,   0.007526,    0.007526,    0.007526,
  0.007503,   0.007503,    0.007503,    0.007503,
  0.007466,   0.007466,    0.007466,    0.007466,
  0.007461,   0.007461,    0.007461,    0.007461,
  0.007461,   0.007461,    0.007461,    0.007461,
  0.007475,   0.007475,    0.007475,    0.007475,
  0.007432,   0.007432,    0.007432,    0.007432,
  0.007311,   0.007311,    0.007311,    0.007311,
  0.007264,   0.007264,    0.007264,    0.007264,
  0.007163,   0.007163,    0.007163,    0.007163,
  0.006826,   0.006826,    0.006826,    0.006826,
  0.00662,    0.00662,     0.00662,     0.00662,
  0.006652,   0.006652,    0.006652,    0.006652,
  0.006567,   0.006567,    0.006567,    0.006567,
  0.006406,   0.006406,    0.006406,    0.006406,
  0.006284,   0.006284,    0.006284,    0.006284,
  0.005968,   0.005968,    0.005968,    0.005968,
  0.005751,   0.005751,    0.005751,    0.005751,
  0.005677,   0.005677,    0.005677,    0.005677,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005589,   0.005589,    0.005589,    0.005589,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005423,   0.005423,    0.005423,    0.005423,
  0.005226,   0.005226,    0.005226,    0.005226,
  0.005117,   0.005117,    0.005117,    0.005117,
  0.005157,   0.005157,    0.005157,    0.005157,
  0.005135,   0.005135,    0.005135,    0.005135,
  0.005079,   0.005079,    0.005079,    0.005079,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005133,   0.005133,    0.005133,    0.005133,
  0.005007,   0.005007,    0.005007,    0.005007,
  0.005082,   0.005082,    0.005082,    0.005082,
  0.005428,   0.005428,    0.005428,    0.005428,
  0.005666,   0.005666,    0.005666,    0.005666,
  0.005685,   0.005685,    0.005685,    0.005685,
  0.005693,   0.005693,    0.005693,    0.005693,
  0.005754,   0.005754,    0.005754,    0.005754,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005874,   0.005874,    0.005874,    0.005874,
  0.005855,   0.005855,    0.005855,    0.005855,
  0.005917,   0.005917,    0.005917,    0.005917,
  0.005963,   0.005963,    0.005963,    0.005963,
  0.005939,   0.005939,    0.005939,    0.005939,
  0.005994,   0.005994,    0.005994,    0.005994,
  0.006069,   0.006069,    0.006069,    0.006069,
  0.006057,   0.006057,    0.006057,    0.006057,
  0.005994,   0.005994,    0.005994,    0.005994,
  0.005954,   0.005954,    0.005954,    0.005954,
  0.006041,   0.006041,    0.006041,    0.006041,
  0.006089,   0.006089,    0.006089,    0.006089,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006172,   0.006172,    0.006172,    0.006172,
  0.006277,   0.006277,    0.006277,    0.006277,
  0.005938,   0.005938,    0.005938,    0.005938,
  0.005406,   0.005406,    0.005406,    0.005406,
  0.00529,    0.00529,     0.00529,     0.00529,
  0.005419,   0.005419,    0.005419,    0.005419,
  0.005482,   0.005482,    0.005482,    0.005482,
  0.005367,   0.005367,    0.005367,    0.005367,
  0.005096,   0.005096,    0.005096,    0.005096,
  0.004927,   0.004927,    0.004927,    0.004927,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004735,   0.004735,    0.004735,    0.004735,
  0.004675,   0.004675,    0.004675,    0.004675,
  0.004672,   0.004672,    0.004672,    0.004672,
  0.00472,    0.00472,     0.00472,     0.00472,
  0.004895,   0.004895,    0.004895,    0.004895,
  0.005025,   0.005025,    0.005025,    0.005025,
  0.005057,   0.005057,    0.005057,    0.005057,
  0.005028,   0.005028,    0.005028,    0.005028,
  0.004963,   0.004963,    0.004963,    0.004963,
  0.005015,   0.005015,    0.005015,    0.005015,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005147,   0.005147,    0.005147,    0.005147,
  0.005157,   0.005157,    0.005157,    0.005157,
  0.005159,   0.005159,    0.005159,    0.005159,
  0.005196,   0.005196,    0.005196,    0.005196,
  0.005274,   0.005274,    0.005274,    0.005274,
  0.005393,   0.005393,    0.005393,    0.005393,
  0.005537,   0.005537,    0.005537,    0.005537,
  0.005743,   0.005743,    0.005743,    0.005743,
  0.005906,   0.005906,    0.005906,    0.005906,
  0.005918,   0.005918,    0.005918,    0.005918,
  0.005932,   0.005932,    0.005932,    0.005932,
  0.005988,   0.005988,    0.005988,    0.005988,
  0.00598,    0.00598,     0.00598,     0.00598,
  0.005916,   0.005916,    0.005916,    0.005916,
  0.005857,   0.005857,    0.005857,    0.005857,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005848,   0.005848,    0.005848,    0.005848,
  0.005782,   0.005782,    0.005782,    0.005782,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005623,   0.005623,    0.005623,    0.005623,
  0.005587,   0.005587,    0.005587,    0.005587,
  0.005573,   0.005573,    0.005573,    0.005573,
  0.00555,    0.00555,     0.00555,     0.00555,
  0.005555,   0.005555,    0.005555,    0.005555,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005631,   0.005631,    0.005631,    0.005631,
  0.005814,   0.005814,    0.005814,    0.005814,
  0.005951,   0.005951,    0.005951,    0.005951,
  0.005992,   0.005992,    0.005992,    0.005992,
  0.006016,   0.006016,    0.006016,    0.006016,
  0.005901,   0.005901,    0.005901,    0.005901,
  0.005676,   0.005676,    0.005676,    0.005676,
  0.005517,   0.005517,    0.005517,    0.005517,
  0.005459,   0.005459,    0.005459,    0.005459,
  0.005384,   0.005384,    0.005384,    0.005384,
  0.005348,   0.005348,    0.005348,    0.005348,
  0.005284,   0.005284,    0.005284,    0.005284,
  0.005072,   0.005072,    0.005072,    0.005072,
  0.004939,   0.004939,    0.004939,    0.004939,
  0.004951,   0.004951,    0.004951,    0.004951,
  0.004871,   0.004871,    0.004871,    0.004871,
  0.004789,   0.004789,    0.004789,    0.004789,
  0.004837,   0.004837,    0.004837,    0.004837,
  0.004866,   0.004866,    0.004866,    0.004866,
  0.004801,   0.004801,    0.004801,    0.004801,
  0.00467,    0.00467,     0.00467,     0.00467,
  0.004582,   0.004582,    0.004582,    0.004582,
  0.004517,   0.004517,    0.004517,    0.004517,
  0.004473,   0.004473,    0.004473,    0.004473,
  0.004629,   0.004629,    0.004629,    0.004629,
  0.004938,   0.004938,    0.004938,    0.004938,
  0.005102,   0.005102,    0.005102,    0.005102,
  0.005046,   0.005046,    0.005046,    0.005046,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005155,   0.005155,    0.005155,    0.005155,
  0.00531,    0.00531,     0.00531,     0.00531,
  0.005597,   0.005597,    0.005597,    0.005597,
  0.005672,   0.005672,    0.005672,    0.005672,
  0.005569,   0.005569,    0.005569,    0.005569,
  0.005571,   0.005571,    0.005571,    0.005571,
  0.005636,   0.005636,    0.005636,    0.005636,
  0.005735,   0.005735,    0.005735,    0.005735,
  0.005779,   0.005779,    0.005779,    0.005779,
  0.005748,   0.005748,    0.005748,    0.005748,
  0.00573,    0.00573,     0.00573,     0.00573,
  0.005669,   0.005669,    0.005669,    0.005669,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005659,   0.005659,    0.005659,    0.005659,
  0.005541,   0.005541,    0.005541,    0.005541,
  0.005373,   0.005373,    0.005373,    0.005373,
  0.005401,   0.005401,    0.005401,    0.005401,
  0.005505,   0.005505,    0.005505,    0.005505,
  0.005539,   0.005539,    0.005539,    0.005539,
  0.005571,   0.005571,    0.005571,    0.005571,
  0.005637,   0.005637,    0.005637,    0.005637,
  0.005746,   0.005746,    0.005746,    0.005746,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.006011,   0.006011,    0.006011,    0.006011,
  0.006145,   0.006145,    0.006145,    0.006145,
  0.005805,   0.005805,    0.005805,    0.005805,
  0.005485,   0.005485,    0.005485,    0.005485,
  0.00537,    0.00537,     0.00537,     0.00537,
  0.005471,   0.005471,    0.005471,    0.005471,
  0.005451,   0.005451,    0.005451,    0.005451,
  0.00524,    0.00524,     0.00524,     0.00524,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005131,   0.005131,    0.005131,    0.005131,
  0.004935,   0.004935,    0.004935,    0.004935,
  0.004692,   0.004692,    0.004692,    0.004692,
  0.004524,   0.004524,    0.004524,    0.004524,
  0.004381,   0.004381,    0.004381,    0.004381,
  0.004259,   0.004259,    0.004259,    0.004259,
  0.004211,   0.004211,    0.004211,    0.004211,
  0.004275,   0.004275,    0.004275,    0.004275,
  0.004468,   0.004468,    0.004468,    0.004468,
  0.004429,   0.004429,    0.004429,    0.004429,
  0.004364,   0.004364,    0.004364,    0.004364,
  0.004364,   0.004364,    0.004364,    0.004364,
  0.004365,   0.004365,    0.004365,    0.004365,
  0.004366,   0.004366,    0.004366,    0.004366,
  0.004439,   0.004439,    0.004439,    0.004439,
  0.004456,   0.004456,    0.004456,    0.004456,
  0.004855,   0.004855,    0.004855,    0.004855,
  0.005524,   0.005524,    0.005524,    0.005524,
  0.005778,   0.005778,    0.005778,    0.005778,
  0.005871,   0.005871,    0.005871,    0.005871,
  0.005881,   0.005881,    0.005881,    0.005881,
  0.005914,   0.005914,    0.005914,    0.005914,
  0.005966,   0.005966,    0.005966,    0.005966,
  0.005972,   0.005972,    0.005972,    0.005972,
  0.005961,   0.005961,    0.005961,    0.005961,
  0.005949,   0.005949,    0.005949,    0.005949,
  0.005927,   0.005927,    0.005927,    0.005927,
  0.005895,   0.005895,    0.005895,    0.005895,
  0.005873,   0.005873,    0.005873,    0.005873,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005833,   0.005833,    0.005833,    0.005833,
  0.005836,   0.005836,    0.005836,    0.005836,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.00583,    0.00583,     0.00583,     0.00583,
  0.005802,   0.005802,    0.005802,    0.005802,
  0.005876,   0.005876,    0.005876,    0.005876,
  0.005868,   0.005868,    0.005868,    0.005868,
  0.005656,   0.005656,    0.005656,    0.005656,
  0.005282,   0.005282,    0.005282,    0.005282,
  0.004906,   0.004906,    0.004906,    0.004906,
  0.004665,   0.004665,    0.004665,    0.004665,
  0.00448,    0.00448,     0.00448,     0.00448,
  0.00421,    0.00421,     0.00421,     0.00421,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.003569,   0.003569,    0.003569,    0.003569,
  0.003352,   0.003352,    0.003352,    0.003352,
  0.003293,   0.003293,    0.003293,    0.003293,
  0.003264,   0.003264,    0.003264,    0.003264,
  0.003303,   0.003303,    0.003303,    0.003303,
  0.003343,   0.003343,    0.003343,    0.003343,
  0.003316,   0.003316,    0.003316,    0.003316,
  0.003265,   0.003265,    0.003265,    0.003265,
  0.003128,   0.003128,    0.003128,    0.003128,
  0.003106,   0.003106,    0.003106,    0.003106,
  0.003194,   0.003194,    0.003194,    0.003194,
  0.003226,   0.003226,    0.003226,    0.003226,
  0.003355,   0.003355,    0.003355,    0.003355,
  0.003351,   0.003351,    0.003351,    0.003351,
  0.003411,   0.003411,    0.003411,    0.003411,
  0.003749,   0.003749,    0.003749,    0.003749,
  0.004052,   0.004052,    0.004052,    0.004052,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004438,   0.004438,    0.004438,    0.004438,
  0.004805,   0.004805,    0.004805,    0.004805,
  0.005239,   0.005239,    0.005239,    0.005239,
  0.005528,   0.005528,    0.005528,    0.005528,
  0.005665,   0.005665,    0.005665,    0.005665,
  0.005962,   0.005962,    0.005962,    0.005962,
  0.006558,   0.006558,    0.006558,    0.006558,
  0.007209,   0.007209,    0.007209,    0.007209,
  0.007611,   0.007611,    0.007611,    0.007611,
  0.007777,   0.007777,    0.007777,    0.007777,
  0.007874,   0.007874,    0.007874,    0.007874,
  0.007979,   0.007979,    0.007979,    0.007979,
  0.008094,   0.008094,    0.008094,    0.008094,
  0.008181,   0.008181,    0.008181,    0.008181,
  0.008201,   0.008201,    0.008201,    0.008201,
  0.008122,   0.008122,    0.008122,    0.008122,
  0.007882,   0.007882,    0.007882,    0.007882,
  0.007699,   0.007699,    0.007699,    0.007699,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007575,   0.007575,    0.007575,    0.007575,
  0.007368,   0.007368,    0.007368,    0.007368,
  0.007325,   0.007325,    0.007325,    0.007325,
  0.007378,   0.007378,    0.007378,    0.007378,
  0.007443,   0.007443,    0.007443,    0.007443,
  0.007642,   0.007642,    0.007642,    0.007642,
  0.007859,   0.007859,    0.007859,    0.007859,
  0.007989,   0.007989,    0.007989,    0.007989,
  0.007986,   0.007986,    0.007986,    0.007986,
  0.007786,   0.007786,    0.007786,    0.007786,
  0.007438,   0.007438,    0.007438,    0.007438,
  0.007125,   0.007125,    0.007125,    0.007125,
  0.006869,   0.006869,    0.006869,    0.006869,
  0.006489,   0.006489,    0.006489,    0.006489,
  0.006119,   0.006119,    0.006119,    0.006119,
  0.005831,   0.005831,    0.005831,    0.005831,
  0.005604,   0.005604,    0.005604,    0.005604,
  0.00555,    0.00555,     0.00555,     0.00555,
  0.005523,   0.005523,    0.005523,    0.005523,
  0.005443,   0.005443,    0.005443,    0.005443,
  0.005279,   0.005279,    0.005279,    0.005279,
  0.005252,   0.005252,    0.005252,    0.005252,
  0.005285,   0.005285,    0.005285,    0.005285,
  0.005005,   0.005005,    0.005005,    0.005005,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.00575,    0.00575,     0.00575,     0.00575,
  0.00599,    0.00599,     0.00599,     0.00599,
  0.005858,   0.005858,    0.005858,    0.005858,
  0.005826,   0.005826,    0.005826,    0.005826,
  0.00601,    0.00601,     0.00601,     0.00601,
  0.006348,   0.006348,    0.006348,    0.006348,
  0.006779,   0.006779,    0.006779,    0.006779,
  0.006895,   0.006895,    0.006895,    0.006895,
  0.006974,   0.006974,    0.006974,    0.006974,
  0.007117,   0.007117,    0.007117,    0.007117,
  0.007134,   0.007134,    0.007134,    0.007134,
  0.007137,   0.007137,    0.007137,    0.007137,
  0.007372,   0.007372,    0.007372,    0.007372,
  0.007591,   0.007591,    0.007591,    0.007591,
  0.007645,   0.007645,    0.007645,    0.007645,
  0.007816,   0.007816,    0.007816,    0.007816,
  0.00792,    0.00792,     0.00792,     0.00792,
  0.008159,   0.008159,    0.008159,    0.008159,
  0.008452,   0.008452,    0.008452,    0.008452,
  0.008541,   0.008541,    0.008541,    0.008541,
  0.008597,   0.008597,    0.008597,    0.008597,
  0.008579,   0.008579,    0.008579,    0.008579,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.008629,   0.008629,    0.008629,    0.008629,
  0.008754,   0.008754,    0.008754,    0.008754,
  0.008829,   0.008829,    0.008829,    0.008829,
  0.008797,   0.008797,    0.008797,    0.008797,
  0.008811,   0.008811,    0.008811,    0.008811,
  0.008844,   0.008844,    0.008844,    0.008844,
  0.008699,   0.008699,    0.008699,    0.008699,
  0.008573,   0.008573,    0.008573,    0.008573,
  0.008497,   0.008497,    0.008497,    0.008497,
  0.008236,   0.008236,    0.008236,    0.008236,
  0.007902,   0.007902,    0.007902,    0.007902,
  0.00754,    0.00754,     0.00754,     0.00754,
  0.007131,   0.007131,    0.007131,    0.007131,
  0.006571,   0.006571,    0.006571,    0.006571,
  0.006325,   0.006325,    0.006325,    0.006325,
  0.006772,   0.006772,    0.006772,    0.006772,
  0.007359,   0.007359,    0.007359,    0.007359,
  0.007377,   0.007377,    0.007377,    0.007377,
  0.006918,   0.006918,    0.006918,    0.006918,
  0.006713,   0.006713,    0.006713,    0.006713,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.006473,   0.006473,    0.006473,    0.006473,
  0.006576,   0.006576,    0.006576,    0.006576,
  0.006491,   0.006491,    0.006491,    0.006491,
  0.006522,   0.006522,    0.006522,    0.006522,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006212,   0.006212,    0.006212,    0.006212,
  0.006426,   0.006426,    0.006426,    0.006426,
  0.006814,   0.006814,    0.006814,    0.006814,
  0.0069,     0.0069,      0.0069,      0.0069,
  0.006598,   0.006598,    0.006598,    0.006598,
  0.006479,   0.006479,    0.006479,    0.006479,
  0.006837,   0.006837,    0.006837,    0.006837,
  0.007106,   0.007106,    0.007106,    0.007106,
  0.00713,    0.00713,     0.00713,     0.00713,
  0.007148,   0.007148,    0.007148,    0.007148,
  0.007211,   0.007211,    0.007211,    0.007211,
  0.007266,   0.007266,    0.007266,    0.007266,
  0.00722,    0.00722,     0.00722,     0.00722,
  0.00712,    0.00712,     0.00712,     0.00712,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007182,   0.007182,    0.007182,    0.007182,
  0.007232,   0.007232,    0.007232,    0.007232,
  0.007268,   0.007268,    0.007268,    0.007268,
  0.007191,   0.007191,    0.007191,    0.007191,
  0.007093,   0.007093,    0.007093,    0.007093,
  0.007071,   0.007071,    0.007071,    0.007071,
  0.007099,   0.007099,    0.007099,    0.007099,
  0.00714,    0.00714,     0.00714,     0.00714,
  0.00714,    0.00714,     0.00714,     0.00714,
  0.007147,   0.007147,    0.007147,    0.007147,
  0.007114,   0.007114,    0.007114,    0.007114,
  0.007039,   0.007039,    0.007039,    0.007039,
  0.006949,   0.006949,    0.006949,    0.006949,
  0.006812,   0.006812,    0.006812,    0.006812,
  0.006594,   0.006594,    0.006594,    0.006594,
  0.006282,   0.006282,    0.006282,    0.006282,
  0.006003,   0.006003,    0.006003,    0.006003,
  0.00581,    0.00581,     0.00581,     0.00581,
  0.005796,   0.005796,    0.005796,    0.005796,
  0.005926,   0.005926,    0.005926,    0.005926,
  0.006003,   0.006003,    0.006003,    0.006003,
  0.005992,   0.005992,    0.005992,    0.005992,
  0.006064,   0.006064,    0.006064,    0.006064,
  0.006633,   0.006633,    0.006633,    0.006633,
  0.006866,   0.006866,    0.006866,    0.006866,
  0.006571,   0.006571,    0.006571,    0.006571,
  0.006392,   0.006392,    0.006392,    0.006392,
  0.006199,   0.006199,    0.006199,    0.006199,
  0.006247,   0.006247,    0.006247,    0.006247,
  0.00667,    0.00667,     0.00667,     0.00667,
  0.007332,   0.007332,    0.007332,    0.007332,
  0.00775,    0.00775,     0.00775,     0.00775,
  0.007743,   0.007743,    0.007743,    0.007743,
  0.007679,   0.007679,    0.007679,    0.007679,
  0.007638,   0.007638,    0.007638,    0.007638,
  0.007646,   0.007646,    0.007646,    0.007646,
  0.007559,   0.007559,    0.007559,    0.007559,
  0.007224,   0.007224,    0.007224,    0.007224,
  0.006972,   0.006972,    0.006972,    0.006972,
  0.007006,   0.007006,    0.007006,    0.007006,
  0.007277,   0.007277,    0.007277,    0.007277,
  0.007564,   0.007564,    0.007564,    0.007564,
  0.007591,   0.007591,    0.007591,    0.007591,
  0.007502,   0.007502,    0.007502,    0.007502,
  0.007521,   0.007521,    0.007521,    0.007521,
  0.007575,   0.007575,    0.007575,    0.007575,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007553,   0.007553,    0.007553,    0.007553,
  0.007553,   0.007553,    0.007553,    0.007553,
  0.007553,   0.007553,    0.007553,    0.007553,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007597,   0.007597,    0.007597,    0.007597,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007799,   0.007799,    0.007799,    0.007799,
  0.007936,   0.007936,    0.007936,    0.007936,
  0.008099,   0.008099,    0.008099,    0.008099,
  0.008131,   0.008131,    0.008131,    0.008131,
  0.008047,   0.008047,    0.008047,    0.008047,
  0.007785,   0.007785,    0.007785,    0.007785,
  0.00761,    0.00761,     0.00761,     0.00761,
  0.00784,    0.00784,     0.00784,     0.00784,
  0.007996,   0.007996,    0.007996,    0.007996,
  0.008043,   0.008043,    0.008043,    0.008043,
  0.008114,   0.008114,    0.008114,    0.008114,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008122,   0.008122,    0.008122,    0.008122,
  0.008153,   0.008153,    0.008153,    0.008153,
  0.008106,   0.008106,    0.008106,    0.008106,
  0.008106,   0.008106,    0.008106,    0.008106,
  0.008114,   0.008114,    0.008114,    0.008114,
  0.007988,   0.007988,    0.007988,    0.007988,
  0.007846,   0.007846,    0.007846,    0.007846,
  0.007783,   0.007783,    0.007783,    0.007783,
  0.007705,   0.007705,    0.007705,    0.007705,
  0.007602,   0.007602,    0.007602,    0.007602,
  0.007484,   0.007484,    0.007484,    0.007484,
  0.007343,   0.007343,    0.007343,    0.007343,
  0.007438,   0.007438,    0.007438,    0.007438,
  0.007636,   0.007636,    0.007636,    0.007636,
  0.007629,   0.007629,    0.007629,    0.007629,
  0.007583,   0.007583,    0.007583,    0.007583,
  0.007596,   0.007596,    0.007596,    0.007596,
  0.007632,   0.007632,    0.007632,    0.007632,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007597,   0.007597,    0.007597,    0.007597,
  0.007597,   0.007597,    0.007597,    0.007597,
  0.007597,   0.007597,    0.007597,    0.007597,
  0.007575,   0.007575,    0.007575,    0.007575,
  0.007553,   0.007553,    0.007553,    0.007553,
  0.007531,   0.007531,    0.007531,    0.007531,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.007465,   0.007465,    0.007465,    0.007465,
  0.007433,   0.007433,    0.007433,    0.007433,
  0.007433,   0.007433,    0.007433,    0.007433,
  0.007443,   0.007443,    0.007443,    0.007443,
  0.007421,   0.007421,    0.007421,    0.007421,
  0.00739,    0.00739,     0.00739,     0.00739,
  0.007337,   0.007337,    0.007337,    0.007337,
  0.007293,   0.007293,    0.007293,    0.007293,
  0.007284,   0.007284,    0.007284,    0.007284,
  0.007276,   0.007276,    0.007276,    0.007276,
  0.007247,   0.007247,    0.007247,    0.007247,
  0.007184,   0.007184,    0.007184,    0.007184,
  0.007116,   0.007116,    0.007116,    0.007116,
  0.007003,   0.007003,    0.007003,    0.007003,
  0.006848,   0.006848,    0.006848,    0.006848,
  0.006634,   0.006634,    0.006634,    0.006634,
  0.00632,    0.00632,     0.00632,     0.00632,
  0.006063,   0.006063,    0.006063,    0.006063,
  0.005909,   0.005909,    0.005909,    0.005909,
  0.005875,   0.005875,    0.005875,    0.005875,
  0.005882,   0.005882,    0.005882,    0.005882,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005605,   0.005605,    0.005605,    0.005605,
  0.005643,   0.005643,    0.005643,    0.005643,
  0.005517,   0.005517,    0.005517,    0.005517,
  0.005315,   0.005315,    0.005315,    0.005315,
  0.005263,   0.005263,    0.005263,    0.005263,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.00531,    0.00531,     0.00531,     0.00531,
  0.00527,    0.00527,     0.00527,     0.00527,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005409,   0.005409,    0.005409,    0.005409,
  0.005409,   0.005409,    0.005409,    0.005409,
  0.005531,   0.005531,    0.005531,    0.005531,
  0.005573,   0.005573,    0.005573,    0.005573,
  0.005657,   0.005657,    0.005657,    0.005657,
  0.005728,   0.005728,    0.005728,    0.005728,
  0.005752,   0.005752,    0.005752,    0.005752,
  0.005659,   0.005659,    0.005659,    0.005659,
  0.005531,   0.005531,    0.005531,    0.005531,
  0.005569,   0.005569,    0.005569,    0.005569,
  0.005603,   0.005603,    0.005603,    0.005603,
  0.005622,   0.005622,    0.005622,    0.005622,
  0.005663,   0.005663,    0.005663,    0.005663,
  0.005713,   0.005713,    0.005713,    0.005713,
  0.005739,   0.005739,    0.005739,    0.005739,
  0.00571,    0.00571,     0.00571,     0.00571,
  0.005666,   0.005666,    0.005666,    0.005666,
  0.005667,   0.005667,    0.005667,    0.005667,
  0.005677,   0.005677,    0.005677,    0.005677,
  0.005699,   0.005699,    0.005699,    0.005699,
  0.005677,   0.005677,    0.005677,    0.005677,
  0.005581,   0.005581,    0.005581,    0.005581,
  0.005436,   0.005436,    0.005436,    0.005436,
  0.005331,   0.005331,    0.005331,    0.005331,
  0.005381,   0.005381,    0.005381,    0.005381,
  0.005464,   0.005464,    0.005464,    0.005464,
  0.00558,    0.00558,     0.00558,     0.00558,
  0.005824,   0.005824,    0.005824,    0.005824,
  0.00613,    0.00613,     0.00613,     0.00613,
  0.006224,   0.006224,    0.006224,    0.006224,
  0.005982,   0.005982,    0.005982,    0.005982,
  0.005755,   0.005755,    0.005755,    0.005755,
  0.005434,   0.005434,    0.005434,    0.005434,
  0.005145,   0.005145,    0.005145,    0.005145,
  0.005195,   0.005195,    0.005195,    0.005195,
  0.005231,   0.005231,    0.005231,    0.005231,
  0.005061,   0.005061,    0.005061,    0.005061,
  0.00479,    0.00479,     0.00479,     0.00479,
  0.004581,   0.004581,    0.004581,    0.004581,
  0.004598,   0.004598,    0.004598,    0.004598,
  0.004716,   0.004716,    0.004716,    0.004716,
  0.004614,   0.004614,    0.004614,    0.004614,
  0.004548,   0.004548,    0.004548,    0.004548,
  0.004808,   0.004808,    0.004808,    0.004808,
  0.005171,   0.005171,    0.005171,    0.005171,
  0.005434,   0.005434,    0.005434,    0.005434,
  0.005634,   0.005634,    0.005634,    0.005634,
  0.005791,   0.005791,    0.005791,    0.005791,
  0.005921,   0.005921,    0.005921,    0.005921,
  0.006506,   0.006506,    0.006506,    0.006506,
  0.007155,   0.007155,    0.007155,    0.007155,
  0.007492,   0.007492,    0.007492,    0.007492,
  0.007808,   0.007808,    0.007808,    0.007808,
  0.007949,   0.007949,    0.007949,    0.007949,
  0.007957,   0.007957,    0.007957,    0.007957,
  0.007927,   0.007927,    0.007927,    0.007927,
  0.00789,    0.00789,     0.00789,     0.00789,
  0.007799,   0.007799,    0.007799,    0.007799,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007597,   0.007597,    0.007597,    0.007597,
  0.007531,   0.007531,    0.007531,    0.007531,
  0.007531,   0.007531,    0.007531,    0.007531,
  0.007553,   0.007553,    0.007553,    0.007553,
  0.007575,   0.007575,    0.007575,    0.007575,
  0.007641,   0.007641,    0.007641,    0.007641,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007708,   0.007708,    0.007708,    0.007708,
  0.007753,   0.007753,    0.007753,    0.007753,
  0.007776,   0.007776,    0.007776,    0.007776,
  0.007776,   0.007776,    0.007776,    0.007776,
  0.007776,   0.007776,    0.007776,    0.007776,
  0.007799,   0.007799,    0.007799,    0.007799,
  0.007821,   0.007821,    0.007821,    0.007821,
  0.007844,   0.007844,    0.007844,    0.007844,
  0.00789,    0.00789,     0.00789,     0.00789,
  0.007982,   0.007982,    0.007982,    0.007982,
  0.008075,   0.008075,    0.008075,    0.008075,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008145,   0.008145,    0.008145,    0.008145,
  0.008216,   0.008216,    0.008216,    0.008216,
  0.008312,   0.008312,    0.008312,    0.008312,
  0.008457,   0.008457,    0.008457,    0.008457,
  0.008654,   0.008654,    0.008654,    0.008654,
  0.00888,    0.00888,     0.00888,     0.00888,
  0.009056,   0.009056,    0.009056,    0.009056,
  0.009036,   0.009036,    0.009036,    0.009036,
  0.008966,   0.008966,    0.008966,    0.008966,
  0.009012,   0.009012,    0.009012,    0.009012,
  0.009059,   0.009059,    0.009059,    0.009059,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.009137,   0.009137,    0.009137,    0.009137,
  0.009147,   0.009147,    0.009147,    0.009147,
  0.00919,    0.00919,     0.00919,     0.00919,
  0.009383,   0.009383,    0.009383,    0.009383,
  0.009342,   0.009342,    0.009342,    0.009342,
  0.009149,   0.009149,    0.009149,    0.009149,
  0.009215,   0.009215,    0.009215,    0.009215,
  0.009345,   0.009345,    0.009345,    0.009345,
  0.009194,   0.009194,    0.009194,    0.009194,
  0.008991,   0.008991,    0.008991,    0.008991,
  0.008943,   0.008943,    0.008943,    0.008943,
  0.00886,    0.00886,     0.00886,     0.00886,
  0.008773,   0.008773,    0.008773,    0.008773,
  0.008678,   0.008678,    0.008678,    0.008678,
  0.008584,   0.008584,    0.008584,    0.008584,
  0.008572,   0.008572,    0.008572,    0.008572,
  0.008506,   0.008506,    0.008506,    0.008506,
  0.008384,   0.008384,    0.008384,    0.008384,
  0.008336,   0.008336,    0.008336,    0.008336,
  0.00836,    0.00836,     0.00836,     0.00836,
  0.008408,   0.008408,    0.008408,    0.008408,
  0.008432,   0.008432,    0.008432,    0.008432,
  0.008432,   0.008432,    0.008432,    0.008432,
  0.008457,   0.008457,    0.008457,    0.008457,
  0.008481,   0.008481,    0.008481,    0.008481,
  0.008506,   0.008506,    0.008506,    0.008506,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.008629,   0.008629,    0.008629,    0.008629,
  0.008754,   0.008754,    0.008754,    0.008754,
  0.00888,    0.00888,     0.00888,     0.00888,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.009216,   0.009216,    0.009216,    0.009216,
  0.00928,    0.00928,     0.00928,     0.00928,
  0.009212,   0.009212,    0.009212,    0.009212,
  0.009003,   0.009003,    0.009003,    0.009003,
  0.008706,   0.008706,    0.008706,    0.008706,
  0.008242,   0.008242,    0.008242,    0.008242,
  0.007824,   0.007824,    0.007824,    0.007824,
  0.007418,   0.007418,    0.007418,    0.007418,
  0.007016,   0.007016,    0.007016,    0.007016,
  0.006987,   0.006987,    0.006987,    0.006987,
  0.007268,   0.007268,    0.007268,    0.007268,
  0.007356,   0.007356,    0.007356,    0.007356,
  0.007462,   0.007462,    0.007462,    0.007462,
  0.007772,   0.007772,    0.007772,    0.007772,
  0.007848,   0.007848,    0.007848,    0.007848,
  0.007974,   0.007974,    0.007974,    0.007974,
  0.008169,   0.008169,    0.008169,    0.008169,
  0.008249,   0.008249,    0.008249,    0.008249,
  0.008317,   0.008317,    0.008317,    0.008317,
  0.00839,    0.00839,     0.00839,     0.00839,
  0.008513,   0.008513,    0.008513,    0.008513,
  0.008586,   0.008586,    0.008586,    0.008586,
  0.008488,   0.008488,    0.008488,    0.008488,
  0.008377,   0.008377,    0.008377,    0.008377,
  0.008142,   0.008142,    0.008142,    0.008142,
  0.007786,   0.007786,    0.007786,    0.007786,
  0.007515,   0.007515,    0.007515,    0.007515,
  0.007327,   0.007327,    0.007327,    0.007327,
  0.007257,   0.007257,    0.007257,    0.007257,
  0.007317,   0.007317,    0.007317,    0.007317,
  0.007358,   0.007358,    0.007358,    0.007358,
  0.007358,   0.007358,    0.007358,    0.007358,
  0.007305,   0.007305,    0.007305,    0.007305,
  0.007166,   0.007166,    0.007166,    0.007166,
  0.00705,    0.00705,     0.00705,     0.00705,
  0.007124,   0.007124,    0.007124,    0.007124,
  0.007315,   0.007315,    0.007315,    0.007315,
  0.007414,   0.007414,    0.007414,    0.007414,
  0.007436,   0.007436,    0.007436,    0.007436,
  0.007424,   0.007424,    0.007424,    0.007424,
  0.007433,   0.007433,    0.007433,    0.007433,
  0.007531,   0.007531,    0.007531,    0.007531,
  0.007637,   0.007637,    0.007637,    0.007637,
  0.007684,   0.007684,    0.007684,    0.007684,
  0.007729,   0.007729,    0.007729,    0.007729,
  0.007814,   0.007814,    0.007814,    0.007814,
  0.007879,   0.007879,    0.007879,    0.007879,
  0.007874,   0.007874,    0.007874,    0.007874,
  0.007789,   0.007789,    0.007789,    0.007789,
  0.007733,   0.007733,    0.007733,    0.007733,
  0.007798,   0.007798,    0.007798,    0.007798,
  0.007932,   0.007932,    0.007932,    0.007932,
  0.008054,   0.008054,    0.008054,    0.008054,
  0.008088,   0.008088,    0.008088,    0.008088,
  0.007874,   0.007874,    0.007874,    0.007874,
  0.007744,   0.007744,    0.007744,    0.007744,
  0.008143,   0.008143,    0.008143,    0.008143,
  0.008475,   0.008475,    0.008475,    0.008475,
  0.008683,   0.008683,    0.008683,    0.008683,
  0.008576,   0.008576,    0.008576,    0.008576,
  0.008454,   0.008454,    0.008454,    0.008454,
  0.008667,   0.008667,    0.008667,    0.008667,
  0.008434,   0.008434,    0.008434,    0.008434,
  0.008218,   0.008218,    0.008218,    0.008218,
  0.008212,   0.008212,    0.008212,    0.008212,
  0.008167,   0.008167,    0.008167,    0.008167,
  0.008261,   0.008261,    0.008261,    0.008261,
  0.008043,   0.008043,    0.008043,    0.008043,
  0.007424,   0.007424,    0.007424,    0.007424,
  0.007049,   0.007049,    0.007049,    0.007049,
  0.007135,   0.007135,    0.007135,    0.007135,
  0.007161,   0.007161,    0.007161,    0.007161,
  0.007034,   0.007034,    0.007034,    0.007034,
  0.007077,   0.007077,    0.007077,    0.007077,
  0.007239,   0.007239,    0.007239,    0.007239,
  0.007386,   0.007386,    0.007386,    0.007386,
  0.007331,   0.007331,    0.007331,    0.007331,
  0.007243,   0.007243,    0.007243,    0.007243,
  0.007182,   0.007182,    0.007182,    0.007182,
  0.007048,   0.007048,    0.007048,    0.007048,
  0.006928,   0.006928,    0.006928,    0.006928,
  0.006856,   0.006856,    0.006856,    0.006856,
  0.00676,    0.00676,     0.00676,     0.00676,
  0.006723,   0.006723,    0.006723,    0.006723,
  0.006733,   0.006733,    0.006733,    0.006733,
  0.00677,    0.00677,     0.00677,     0.00677,
  0.006863,   0.006863,    0.006863,    0.006863,
  0.006941,   0.006941,    0.006941,    0.006941,
  0.007012,   0.007012,    0.007012,    0.007012,
  0.007122,   0.007122,    0.007122,    0.007122,
  0.007284,   0.007284,    0.007284,    0.007284,
  0.007423,   0.007423,    0.007423,    0.007423,
  0.007553,   0.007553,    0.007553,    0.007553,
  0.007736,   0.007736,    0.007736,    0.007736,
  0.007851,   0.007851,    0.007851,    0.007851,
  0.007773,   0.007773,    0.007773,    0.007773,
  0.007678,   0.007678,    0.007678,    0.007678,
  0.007792,   0.007792,    0.007792,    0.007792,
  0.007874,   0.007874,    0.007874,    0.007874,
  0.007737,   0.007737,    0.007737,    0.007737,
  0.007485,   0.007485,    0.007485,    0.007485,
  0.007201,   0.007201,    0.007201,    0.007201,
  0.006903,   0.006903,    0.006903,    0.006903,
  0.006834,   0.006834,    0.006834,    0.006834,
  0.007284,   0.007284,    0.007284,    0.007284,
  0.008504,   0.008504,    0.008504,    0.008504,
  0.009555,   0.009555,    0.009555,    0.009555,
  0.009744,   0.009744,    0.009744,    0.009744,
  0.009792,   0.009792,    0.009792,    0.009792,
  0.009886,   0.009886,    0.009886,    0.009886,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.009942,   0.009942,    0.009942,    0.009942,
  0.009974,   0.009974,    0.009974,    0.009974,
  0.01001,    0.01001,     0.01001,     0.01001,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.009776,   0.009776,    0.009776,    0.009776,
  0.009558,   0.009558,    0.009558,    0.009558,
  0.009562,   0.009562,    0.009562,    0.009562,
  0.009535,   0.009535,    0.009535,    0.009535,
  0.009481,   0.009481,    0.009481,    0.009481,
  0.009454,   0.009454,    0.009454,    0.009454,
  0.009454,   0.009454,    0.009454,    0.009454,
  0.009454,   0.009454,    0.009454,    0.009454,
  0.009454,   0.009454,    0.009454,    0.009454,
  0.009454,   0.009454,    0.009454,    0.009454,
  0.009454,   0.009454,    0.009454,    0.009454,
  0.009428,   0.009428,    0.009428,    0.009428,
  0.009348,   0.009348,    0.009348,    0.009348,
  0.009242,   0.009242,    0.009242,    0.009242,
  0.009137,   0.009137,    0.009137,    0.009137,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.009059,   0.009059,    0.009059,    0.009059,
  0.009033,   0.009033,    0.009033,    0.009033,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.008905,   0.008905,    0.008905,    0.008905,
  0.008905,   0.008905,    0.008905,    0.008905,
  0.008956,   0.008956,    0.008956,    0.008956,
  0.009008,   0.009008,    0.009008,    0.009008,
  0.008991,   0.008991,    0.008991,    0.008991,
  0.008885,   0.008885,    0.008885,    0.008885,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008596,   0.008596,    0.008596,    0.008596,
  0.00858,    0.00858,     0.00858,     0.00858,
  0.008556,   0.008556,    0.008556,    0.008556,
  0.008451,   0.008451,    0.008451,    0.008451,
  0.008398,   0.008398,    0.008398,    0.008398,
  0.008366,   0.008366,    0.008366,    0.008366,
  0.00833,    0.00833,     0.00833,     0.00833,
  0.008325,   0.008325,    0.008325,    0.008325,
  0.008347,   0.008347,    0.008347,    0.008347,
  0.008334,   0.008334,    0.008334,    0.008334,
  0.008307,   0.008307,    0.008307,    0.008307,
  0.008257,   0.008257,    0.008257,    0.008257,
  0.0081,     0.0081,      0.0081,      0.0081,
  0.008001,   0.008001,    0.008001,    0.008001,
  0.008028,   0.008028,    0.008028,    0.008028,
  0.007984,   0.007984,    0.007984,    0.007984,
  0.00795,    0.00795,     0.00795,     0.00795,
  0.008184,   0.008184,    0.008184,    0.008184,
  0.008489,   0.008489,    0.008489,    0.008489,
  0.008542,   0.008542,    0.008542,    0.008542,
  0.008313,   0.008313,    0.008313,    0.008313,
  0.008145,   0.008145,    0.008145,    0.008145,
  0.008169,   0.008169,    0.008169,    0.008169,
  0.008169,   0.008169,    0.008169,    0.008169,
  0.008145,   0.008145,    0.008145,    0.008145,
  0.008145,   0.008145,    0.008145,    0.008145,
  0.008122,   0.008122,    0.008122,    0.008122,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008075,   0.008075,    0.008075,    0.008075,
  0.008005,   0.008005,    0.008005,    0.008005,
  0.007822,   0.007822,    0.007822,    0.007822,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.0074,     0.0074,      0.0074,      0.0074,
  0.007356,   0.007356,    0.007356,    0.007356,
  0.007335,   0.007335,    0.007335,    0.007335,
  0.007356,   0.007356,    0.007356,    0.007356,
  0.00751,    0.00751,     0.00751,     0.00751,
  0.007731,   0.007731,    0.007731,    0.007731,
  0.007844,   0.007844,    0.007844,    0.007844,
  0.007959,   0.007959,    0.007959,    0.007959,
  0.008083,   0.008083,    0.008083,    0.008083,
  0.008091,   0.008091,    0.008091,    0.008091,
  0.008052,   0.008052,    0.008052,    0.008052,
  0.007999,   0.007999,    0.007999,    0.007999,
  0.007851,   0.007851,    0.007851,    0.007851,
  0.007798,   0.007798,    0.007798,    0.007798,
  0.007841,   0.007841,    0.007841,    0.007841,
  0.007817,   0.007817,    0.007817,    0.007817,
  0.007727,   0.007727,    0.007727,    0.007727,
  0.007557,   0.007557,    0.007557,    0.007557,
  0.007328,   0.007328,    0.007328,    0.007328,
  0.007247,   0.007247,    0.007247,    0.007247,
  0.007075,   0.007075,    0.007075,    0.007075,
  0.006375,   0.006375,    0.006375,    0.006375,
  0.005904,   0.005904,    0.005904,    0.005904,
  0.005719,   0.005719,    0.005719,    0.005719,
  0.005565,   0.005565,    0.005565,    0.005565,
  0.005627,   0.005627,    0.005627,    0.005627,
  0.006661,   0.006661,    0.006661,    0.006661,
  0.008108,   0.008108,    0.008108,    0.008108,
  0.008619,   0.008619,    0.008619,    0.008619,
  0.00871,    0.00871,     0.00871,     0.00871,
  0.008806,   0.008806,    0.008806,    0.008806,
  0.008802,   0.008802,    0.008802,    0.008802,
  0.008933,   0.008933,    0.008933,    0.008933,
  0.009044,   0.009044,    0.009044,    0.009044,
  0.00887,    0.00887,     0.00887,     0.00887,
  0.008698,   0.008698,    0.008698,    0.008698,
  0.008446,   0.008446,    0.008446,    0.008446,
  0.008164,   0.008164,    0.008164,    0.008164,
  0.008006,   0.008006,    0.008006,    0.008006,
  0.007901,   0.007901,    0.007901,    0.007901,
  0.007777,   0.007777,    0.007777,    0.007777,
  0.007738,   0.007738,    0.007738,    0.007738,
  0.007715,   0.007715,    0.007715,    0.007715,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007461,   0.007461,    0.007461,    0.007461,
  0.007156,   0.007156,    0.007156,    0.007156,
  0.006998,   0.006998,    0.006998,    0.006998,
  0.006916,   0.006916,    0.006916,    0.006916,
  0.006835,   0.006835,    0.006835,    0.006835,
  0.006795,   0.006795,    0.006795,    0.006795,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006917,   0.006917,    0.006917,    0.006917,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007445,   0.007445,    0.007445,    0.007445,
  0.00787,    0.00787,     0.00787,     0.00787,
  0.008224,   0.008224,    0.008224,    0.008224,
  0.008203,   0.008203,    0.008203,    0.008203,
  0.007986,   0.007986,    0.007986,    0.007986,
  0.007904,   0.007904,    0.007904,    0.007904,
  0.007906,   0.007906,    0.007906,    0.007906,
  0.007866,   0.007866,    0.007866,    0.007866,
  0.007739,   0.007739,    0.007739,    0.007739,
  0.007475,   0.007475,    0.007475,    0.007475,
  0.007097,   0.007097,    0.007097,    0.007097,
  0.006756,   0.006756,    0.006756,    0.006756,
  0.00652,    0.00652,     0.00652,     0.00652,
  0.006349,   0.006349,    0.006349,    0.006349,
  0.006326,   0.006326,    0.006326,    0.006326,
  0.006505,   0.006505,    0.006505,    0.006505,
  0.006461,   0.006461,    0.006461,    0.006461,
  0.006422,   0.006422,    0.006422,    0.006422,
  0.006792,   0.006792,    0.006792,    0.006792,
  0.007261,   0.007261,    0.007261,    0.007261,
  0.007698,   0.007698,    0.007698,    0.007698,
  0.008313,   0.008313,    0.008313,    0.008313,
  0.008991,   0.008991,    0.008991,    0.008991,
  0.009286,   0.009286,    0.009286,    0.009286,
  0.009338,   0.009338,    0.009338,    0.009338,
  0.009428,   0.009428,    0.009428,    0.009428,
  0.009451,   0.009451,    0.009451,    0.009451,
  0.009396,   0.009396,    0.009396,    0.009396,
  0.009378,   0.009378,    0.009378,    0.009378,
  0.009315,   0.009315,    0.009315,    0.009315,
  0.00927,    0.00927,     0.00927,     0.00927,
  0.009258,   0.009258,    0.009258,    0.009258,
  0.009123,   0.009123,    0.009123,    0.009123,
  0.00892,    0.00892,     0.00892,     0.00892,
  0.008716,   0.008716,    0.008716,    0.008716,
  0.008485,   0.008485,    0.008485,    0.008485,
  0.008282,   0.008282,    0.008282,    0.008282,
  0.00813,    0.00813,     0.00813,     0.00813,
  0.007925,   0.007925,    0.007925,    0.007925,
  0.007693,   0.007693,    0.007693,    0.007693,
  0.007538,   0.007538,    0.007538,    0.007538,
  0.007477,   0.007477,    0.007477,    0.007477,
  0.0074,     0.0074,      0.0074,      0.0074,
  0.007292,   0.007292,    0.007292,    0.007292,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007379,   0.007379,    0.007379,    0.007379,
  0.007616,   0.007616,    0.007616,    0.007616,
  0.007761,   0.007761,    0.007761,    0.007761,
  0.007849,   0.007849,    0.007849,    0.007849,
  0.007886,   0.007886,    0.007886,    0.007886,
  0.007806,   0.007806,    0.007806,    0.007806,
  0.007576,   0.007576,    0.007576,    0.007576,
  0.007197,   0.007197,    0.007197,    0.007197,
  0.006872,   0.006872,    0.006872,    0.006872,
  0.006731,   0.006731,    0.006731,    0.006731,
  0.006525,   0.006525,    0.006525,    0.006525,
  0.006445,   0.006445,    0.006445,    0.006445,
  0.006444,   0.006444,    0.006444,    0.006444,
  0.006281,   0.006281,    0.006281,    0.006281,
  0.006025,   0.006025,    0.006025,    0.006025,
  0.005584,   0.005584,    0.005584,    0.005584,
  0.005584,   0.005584,    0.005584,    0.005584,
  0.005931,   0.005931,    0.005931,    0.005931,
  0.005931,   0.005931,    0.005931,    0.005931,
  0.005963,   0.005963,    0.005963,    0.005963,
  0.005806,   0.005806,    0.005806,    0.005806,
  0.005648,   0.005648,    0.005648,    0.005648,
  0.00568,    0.00568,     0.00568,     0.00568,
  0.005649,   0.005649,    0.005649,    0.005649,
  0.0059,     0.0059,      0.0059,      0.0059,
  0.006151,   0.006151,    0.006151,    0.006151,
  0.006404,   0.006404,    0.006404,    0.006404,
  0.006775,   0.006775,    0.006775,    0.006775,
  0.007143,   0.007143,    0.007143,    0.007143,
  0.007364,   0.007364,    0.007364,    0.007364,
  0.007307,   0.007307,    0.007307,    0.007307,
  0.007192,   0.007192,    0.007192,    0.007192,
  0.007169,   0.007169,    0.007169,    0.007169,
  0.007187,   0.007187,    0.007187,    0.007187,
  0.007265,   0.007265,    0.007265,    0.007265,
  0.007374,   0.007374,    0.007374,    0.007374,
  0.007523,   0.007523,    0.007523,    0.007523,
  0.007665,   0.007665,    0.007665,    0.007665,
  0.00772,    0.00772,     0.00772,     0.00772,
  0.007684,   0.007684,    0.007684,    0.007684,
  0.00761,    0.00761,     0.00761,     0.00761,
  0.007507,   0.007507,    0.007507,    0.007507,
  0.007414,   0.007414,    0.007414,    0.007414,
  0.00739,    0.00739,     0.00739,     0.00739,
  0.007292,   0.007292,    0.007292,    0.007292,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007401,   0.007401,    0.007401,    0.007401,
  0.007865,   0.007865,    0.007865,    0.007865,
  0.008188,   0.008188,    0.008188,    0.008188,
  0.008164,   0.008164,    0.008164,    0.008164,
  0.008036,   0.008036,    0.008036,    0.008036,
  0.008043,   0.008043,    0.008043,    0.008043,
  0.00796,    0.00796,     0.00796,     0.00796,
  0.0076,     0.0076,      0.0076,      0.0076,
  0.007293,   0.007293,    0.007293,    0.007293,
  0.006814,   0.006814,    0.006814,    0.006814,
  0.006246,   0.006246,    0.006246,    0.006246,
  0.006089,   0.006089,    0.006089,    0.006089,
  0.006122,   0.006122,    0.006122,    0.006122,
  0.006216,   0.006216,    0.006216,    0.006216,
  0.007136,   0.007136,    0.007136,    0.007136,
  0.007735,   0.007735,    0.007735,    0.007735,
  0.00698,    0.00698,     0.00698,     0.00698,
  0.006246,   0.006246,    0.006246,    0.006246,
  0.005979,   0.005979,    0.005979,    0.005979,
  0.005834,   0.005834,    0.005834,    0.005834,
  0.005742,   0.005742,    0.005742,    0.005742,
  0.005592,   0.005592,    0.005592,    0.005592,
  0.00558,    0.00558,     0.00558,     0.00558,
  0.005927,   0.005927,    0.005927,    0.005927,
  0.006731,   0.006731,    0.006731,    0.006731,
  0.007493,   0.007493,    0.007493,    0.007493,
  0.007921,   0.007921,    0.007921,    0.007921,
  0.00816,    0.00816,     0.00816,     0.00816,
  0.008024,   0.008024,    0.008024,    0.008024,
  0.007983,   0.007983,    0.007983,    0.007983,
  0.008137,   0.008137,    0.008137,    0.008137,
  0.008015,   0.008015,    0.008015,    0.008015,
  0.007688,   0.007688,    0.007688,    0.007688,
  0.007594,   0.007594,    0.007594,    0.007594,
  0.007709,   0.007709,    0.007709,    0.007709,
  0.008025,   0.008025,    0.008025,    0.008025,
  0.008331,   0.008331,    0.008331,    0.008331,
  0.008413,   0.008413,    0.008413,    0.008413,
  0.008338,   0.008338,    0.008338,    0.008338,
  0.008195,   0.008195,    0.008195,    0.008195,
  0.008152,   0.008152,    0.008152,    0.008152,
  0.008114,   0.008114,    0.008114,    0.008114,
  0.008055,   0.008055,    0.008055,    0.008055,
  0.007989,   0.007989,    0.007989,    0.007989,
  0.007934,   0.007934,    0.007934,    0.007934,
  0.007919,   0.007919,    0.007919,    0.007919,
  0.007904,   0.007904,    0.007904,    0.007904,
  0.007919,   0.007919,    0.007919,    0.007919,
  0.007971,   0.007971,    0.007971,    0.007971,
  0.008031,   0.008031,    0.008031,    0.008031,
  0.008119,   0.008119,    0.008119,    0.008119,
  0.008263,   0.008263,    0.008263,    0.008263,
  0.008303,   0.008303,    0.008303,    0.008303,
  0.008224,   0.008224,    0.008224,    0.008224,
  0.008417,   0.008417,    0.008417,    0.008417,
  0.00843,    0.00843,     0.00843,     0.00843,
  0.007888,   0.007888,    0.007888,    0.007888,
  0.007541,   0.007541,    0.007541,    0.007541,
  0.007727,   0.007727,    0.007727,    0.007727,
  0.007827,   0.007827,    0.007827,    0.007827,
  0.007733,   0.007733,    0.007733,    0.007733,
  0.007973,   0.007973,    0.007973,    0.007973,
  0.008279,   0.008279,    0.008279,    0.008279,
  0.008727,   0.008727,    0.008727,    0.008727,
  0.00931,    0.00931,     0.00931,     0.00931,
  0.009571,   0.009571,    0.009571,    0.009571,
  0.009508,   0.009508,    0.009508,    0.009508,
  0.009266,   0.009266,    0.009266,    0.009266,
  0.009041,   0.009041,    0.009041,    0.009041,
  0.009119,   0.009119,    0.009119,    0.009119,
  0.009502,   0.009502,    0.009502,    0.009502,
  0.00961,    0.00961,     0.00961,     0.00961,
  0.009519,   0.009519,    0.009519,    0.009519,
  0.009202,   0.009202,    0.009202,    0.009202,
  0.008649,   0.008649,    0.008649,    0.008649,
  0.008295,   0.008295,    0.008295,    0.008295,
  0.008161,   0.008161,    0.008161,    0.008161,
  0.008116,   0.008116,    0.008116,    0.008116,
  0.008062,   0.008062,    0.008062,    0.008062,
  0.007993,   0.007993,    0.007993,    0.007993,
  0.007939,   0.007939,    0.007939,    0.007939,
  0.00788,    0.00788,     0.00788,     0.00788,
  0.007823,   0.007823,    0.007823,    0.007823,
  0.007723,   0.007723,    0.007723,    0.007723,
  0.007673,   0.007673,    0.007673,    0.007673,
  0.00775,    0.00775,     0.00775,     0.00775,
  0.007764,   0.007764,    0.007764,    0.007764,
  0.007682,   0.007682,    0.007682,    0.007682,
  0.007588,   0.007588,    0.007588,    0.007588,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.007335,   0.007335,    0.007335,    0.007335,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007186,   0.007186,    0.007186,    0.007186,
  0.00725,    0.00725,     0.00725,     0.00725,
  0.007335,   0.007335,    0.007335,    0.007335,
  0.007421,   0.007421,    0.007421,    0.007421,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007624,   0.007624,    0.007624,    0.007624,
  0.007788,   0.007788,    0.007788,    0.007788,
  0.007769,   0.007769,    0.007769,    0.007769,
  0.007374,   0.007374,    0.007374,    0.007374,
  0.007179,   0.007179,    0.007179,    0.007179,
  0.007116,   0.007116,    0.007116,    0.007116,
  0.006888,   0.006888,    0.006888,    0.006888,
  0.006884,   0.006884,    0.006884,    0.006884,
  0.006919,   0.006919,    0.006919,    0.006919,
  0.006821,   0.006821,    0.006821,    0.006821,
  0.006963,   0.006963,    0.006963,    0.006963,
  0.00705,    0.00705,     0.00705,     0.00705,
  0.006967,   0.006967,    0.006967,    0.006967,
  0.00727,    0.00727,     0.00727,     0.00727,
  0.007704,   0.007704,    0.007704,    0.007704,
  0.008073,   0.008073,    0.008073,    0.008073,
  0.008512,   0.008512,    0.008512,    0.008512,
  0.008771,   0.008771,    0.008771,    0.008771,
  0.008805,   0.008805,    0.008805,    0.008805,
  0.008874,   0.008874,    0.008874,    0.008874,
  0.009008,   0.009008,    0.009008,    0.009008,
  0.009132,   0.009132,    0.009132,    0.009132,
  0.009249,   0.009249,    0.009249,    0.009249,
  0.009319,   0.009319,    0.009319,    0.009319,
  0.009374,   0.009374,    0.009374,    0.009374,
  0.009479,   0.009479,    0.009479,    0.009479,
  0.009585,   0.009585,    0.009585,    0.009585,
  0.009637,   0.009637,    0.009637,    0.009637,
  0.009508,   0.009508,    0.009508,    0.009508,
  0.00931,    0.00931,     0.00931,     0.00931,
  0.009167,   0.009167,    0.009167,    0.009167,
  0.009122,   0.009122,    0.009122,    0.009122,
  0.009176,   0.009176,    0.009176,    0.009176,
  0.009207,   0.009207,    0.009207,    0.009207,
  0.009185,   0.009185,    0.009185,    0.009185,
  0.009127,   0.009127,    0.009127,    0.009127,
  0.009043,   0.009043,    0.009043,    0.009043,
  0.009027,   0.009027,    0.009027,    0.009027,
  0.009011,   0.009011,    0.009011,    0.009011,
  0.008965,   0.008965,    0.008965,    0.008965,
  0.008945,   0.008945,    0.008945,    0.008945,
  0.008925,   0.008925,    0.008925,    0.008925,
  0.008905,   0.008905,    0.008905,    0.008905,
  0.00888,    0.00888,     0.00888,     0.00888,
  0.008829,   0.008829,    0.008829,    0.008829,
  0.008753,   0.008753,    0.008753,    0.008753,
  0.008753,   0.008753,    0.008753,    0.008753,
  0.008747,   0.008747,    0.008747,    0.008747,
  0.008684,   0.008684,    0.008684,    0.008684,
  0.008652,   0.008652,    0.008652,    0.008652,
  0.008652,   0.008652,    0.008652,    0.008652,
  0.00879,    0.00879,     0.00879,     0.00879,
  0.008843,   0.008843,    0.008843,    0.008843,
  0.008726,   0.008726,    0.008726,    0.008726,
  0.008753,   0.008753,    0.008753,    0.008753,
  0.008805,   0.008805,    0.008805,    0.008805,
  0.00883,    0.00883,     0.00883,     0.00883,
  0.008812,   0.008812,    0.008812,    0.008812,
  0.008731,   0.008731,    0.008731,    0.008731,
  0.008797,   0.008797,    0.008797,    0.008797,
  0.008907,   0.008907,    0.008907,    0.008907,
  0.009038,   0.009038,    0.009038,    0.009038,
  0.009126,   0.009126,    0.009126,    0.009126,
  0.009069,   0.009069,    0.009069,    0.009069,
  0.009022,   0.009022,    0.009022,    0.009022,
  0.009071,   0.009071,    0.009071,    0.009071,
  0.009232,   0.009232,    0.009232,    0.009232,
  0.00928,    0.00928,     0.00928,     0.00928,
  0.008973,   0.008973,    0.008973,    0.008973,
  0.008622,   0.008622,    0.008622,    0.008622,
  0.008236,   0.008236,    0.008236,    0.008236,
  0.007574,   0.007574,    0.007574,    0.007574,
  0.007261,   0.007261,    0.007261,    0.007261,
  0.007526,   0.007526,    0.007526,    0.007526,
  0.007859,   0.007859,    0.007859,    0.007859,
  0.008137,   0.008137,    0.008137,    0.008137,
  0.008428,   0.008428,    0.008428,    0.008428,
  0.008701,   0.008701,    0.008701,    0.008701,
  0.008954,   0.008954,    0.008954,    0.008954,
  0.009086,   0.009086,    0.009086,    0.009086,
  0.009064,   0.009064,    0.009064,    0.009064,
  0.008996,   0.008996,    0.008996,    0.008996,
  0.008927,   0.008927,    0.008927,    0.008927,
  0.008964,   0.008964,    0.008964,    0.008964,
  0.009043,   0.009043,    0.009043,    0.009043,
  0.009027,   0.009027,    0.009027,    0.009027,
  0.008991,   0.008991,    0.008991,    0.008991,
  0.0089,     0.0089,      0.0089,      0.0089,
  0.008779,   0.008779,    0.008779,    0.008779,
  0.008703,   0.008703,    0.008703,    0.008703,
  0.008653,   0.008653,    0.008653,    0.008653,
  0.008729,   0.008729,    0.008729,    0.008729,
  0.008931,   0.008931,    0.008931,    0.008931,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.009163,   0.009163,    0.009163,    0.009163,
  0.009237,   0.009237,    0.009237,    0.009237,
  0.009172,   0.009172,    0.009172,    0.009172,
  0.008955,   0.008955,    0.008955,    0.008955,
  0.008782,   0.008782,    0.008782,    0.008782,
  0.008637,   0.008637,    0.008637,    0.008637,
  0.0085,     0.0085,      0.0085,      0.0085,
  0.008434,   0.008434,    0.008434,    0.008434,
  0.008437,   0.008437,    0.008437,    0.008437,
  0.008535,   0.008535,    0.008535,    0.008535,
  0.008619,   0.008619,    0.008619,    0.008619,
  0.008547,   0.008547,    0.008547,    0.008547,
  0.008434,   0.008434,    0.008434,    0.008434,
  0.008346,   0.008346,    0.008346,    0.008346,
  0.008301,   0.008301,    0.008301,    0.008301,
  0.008294,   0.008294,    0.008294,    0.008294,
  0.008266,   0.008266,    0.008266,    0.008266,
  0.008213,   0.008213,    0.008213,    0.008213,
  0.008199,   0.008199,    0.008199,    0.008199,
  0.008213,   0.008213,    0.008213,    0.008213,
  0.00815,    0.00815,     0.00815,     0.00815,
  0.007967,   0.007967,    0.007967,    0.007967,
  0.007916,   0.007916,    0.007916,    0.007916,
  0.008028,   0.008028,    0.008028,    0.008028,
  0.008267,   0.008267,    0.008267,    0.008267,
  0.008722,   0.008722,    0.008722,    0.008722,
  0.009012,   0.009012,    0.009012,    0.009012,
  0.009035,   0.009035,    0.009035,    0.009035,
  0.008898,   0.008898,    0.008898,    0.008898,
  0.008661,   0.008661,    0.008661,    0.008661,
  0.008613,   0.008613,    0.008613,    0.008613,
  0.008774,   0.008774,    0.008774,    0.008774,
  0.008951,   0.008951,    0.008951,    0.008951,
  0.009046,   0.009046,    0.009046,    0.009046,
  0.009117,   0.009117,    0.009117,    0.009117,
  0.0091,     0.0091,      0.0091,      0.0091,
  0.008938,   0.008938,    0.008938,    0.008938,
  0.008824,   0.008824,    0.008824,    0.008824,
  0.008793,   0.008793,    0.008793,    0.008793,
  0.008776,   0.008776,    0.008776,    0.008776,
  0.008765,   0.008765,    0.008765,    0.008765,
  0.008754,   0.008754,    0.008754,    0.008754,
  0.008748,   0.008748,    0.008748,    0.008748,
  0.008754,   0.008754,    0.008754,    0.008754,
  0.008676,   0.008676,    0.008676,    0.008676,
  0.008598,   0.008598,    0.008598,    0.008598,
  0.008572,   0.008572,    0.008572,    0.008572,
  0.008572,   0.008572,    0.008572,    0.008572,
  0.008578,   0.008578,    0.008578,    0.008578,
  0.008584,   0.008584,    0.008584,    0.008584,
  0.008635,   0.008635,    0.008635,    0.008635,
  0.008681,   0.008681,    0.008681,    0.008681,
  0.008596,   0.008596,    0.008596,    0.008596,
  0.008493,   0.008493,    0.008493,    0.008493,
  0.008515,   0.008515,    0.008515,    0.008515,
  0.008463,   0.008463,    0.008463,    0.008463,
  0.008378,   0.008378,    0.008378,    0.008378,
  0.008452,   0.008452,    0.008452,    0.008452,
  0.008541,   0.008541,    0.008541,    0.008541,
  0.008472,   0.008472,    0.008472,    0.008472,
  0.008338,   0.008338,    0.008338,    0.008338,
  0.008137,   0.008137,    0.008137,    0.008137,
  0.0079,     0.0079,      0.0079,      0.0079,
  0.007919,   0.007919,    0.007919,    0.007919,
  0.007979,   0.007979,    0.007979,    0.007979,
  0.008104,   0.008104,    0.008104,    0.008104,
  0.008356,   0.008356,    0.008356,    0.008356,
  0.008297,   0.008297,    0.008297,    0.008297,
  0.007988,   0.007988,    0.007988,    0.007988,
  0.007652,   0.007652,    0.007652,    0.007652,
  0.007345,   0.007345,    0.007345,    0.007345,
  0.007159,   0.007159,    0.007159,    0.007159,
  0.007197,   0.007197,    0.007197,    0.007197,
  0.007234,   0.007234,    0.007234,    0.007234,
  0.007286,   0.007286,    0.007286,    0.007286,
  0.007457,   0.007457,    0.007457,    0.007457,
  0.007637,   0.007637,    0.007637,    0.007637,
  0.00776,    0.00776,     0.00776,     0.00776,
  0.007867,   0.007867,    0.007867,    0.007867,
  0.007937,   0.007937,    0.007937,    0.007937,
  0.007965,   0.007965,    0.007965,    0.007965,
  0.007974,   0.007974,    0.007974,    0.007974,
  0.007987,   0.007987,    0.007987,    0.007987,
  0.008,      0.008,       0.008,       0.008,
  0.007983,   0.007983,    0.007983,    0.007983,
  0.007933,   0.007933,    0.007933,    0.007933,
  0.007864,   0.007864,    0.007864,    0.007864,
  0.007804,   0.007804,    0.007804,    0.007804,
  0.007722,   0.007722,    0.007722,    0.007722,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007597,   0.007597,    0.007597,    0.007597,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.007531,   0.007531,    0.007531,    0.007531,
  0.007531,   0.007531,    0.007531,    0.007531,
  0.007688,   0.007688,    0.007688,    0.007688,
  0.008006,   0.008006,    0.008006,    0.008006,
  0.008265,   0.008265,    0.008265,    0.008265,
  0.008432,   0.008432,    0.008432,    0.008432,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.008678,   0.008678,    0.008678,    0.008678,
  0.008804,   0.008804,    0.008804,    0.008804,
  0.008951,   0.008951,    0.008951,    0.008951,
  0.009016,   0.009016,    0.009016,    0.009016,
  0.008719,   0.008719,    0.008719,    0.008719,
  0.008173,   0.008173,    0.008173,    0.008173,
  0.007928,   0.007928,    0.007928,    0.007928,
  0.008005,   0.008005,    0.008005,    0.008005,
  0.008151,   0.008151,    0.008151,    0.008151,
  0.008096,   0.008096,    0.008096,    0.008096,
  0.007894,   0.007894,    0.007894,    0.007894,
  0.007797,   0.007797,    0.007797,    0.007797,
  0.007902,   0.007902,    0.007902,    0.007902,
  0.007783,   0.007783,    0.007783,    0.007783,
  0.007504,   0.007504,    0.007504,    0.007504,
  0.007533,   0.007533,    0.007533,    0.007533,
  0.00734,    0.00734,     0.00734,     0.00734,
  0.007256,   0.007256,    0.007256,    0.007256,
  0.00735,    0.00735,     0.00735,     0.00735,
  0.00713,    0.00713,     0.00713,     0.00713,
  0.006987,   0.006987,    0.006987,    0.006987,
  0.007034,   0.007034,    0.007034,    0.007034,
  0.007105,   0.007105,    0.007105,    0.007105,
  0.007085,   0.007085,    0.007085,    0.007085,
  0.007136,   0.007136,    0.007136,    0.007136,
  0.007385,   0.007385,    0.007385,    0.007385,
  0.0076,     0.0076,      0.0076,      0.0076,
  0.007797,   0.007797,    0.007797,    0.007797,
  0.008015,   0.008015,    0.008015,    0.008015,
  0.008074,   0.008074,    0.008074,    0.008074,
  0.008017,   0.008017,    0.008017,    0.008017,
  0.007998,   0.007998,    0.007998,    0.007998,
  0.008038,   0.008038,    0.008038,    0.008038,
  0.008076,   0.008076,    0.008076,    0.008076,
  0.008095,   0.008095,    0.008095,    0.008095,
  0.008095,   0.008095,    0.008095,    0.008095,
  0.008061,   0.008061,    0.008061,    0.008061,
  0.008015,   0.008015,    0.008015,    0.008015,
  0.00796,    0.00796,     0.00796,     0.00796,
  0.007875,   0.007875,    0.007875,    0.007875,
  0.007795,   0.007795,    0.007795,    0.007795,
  0.007809,   0.007809,    0.007809,    0.007809,
  0.007851,   0.007851,    0.007851,    0.007851,
  0.007887,   0.007887,    0.007887,    0.007887,
  0.007953,   0.007953,    0.007953,    0.007953,
  0.007988,   0.007988,    0.007988,    0.007988,
  0.007965,   0.007965,    0.007965,    0.007965,
  0.007993,   0.007993,    0.007993,    0.007993,
  0.008047,   0.008047,    0.008047,    0.008047,
  0.00801,    0.00801,     0.00801,     0.00801,
  0.007739,   0.007739,    0.007739,    0.007739,
  0.007265,   0.007265,    0.007265,    0.007265,
  0.006733,   0.006733,    0.006733,    0.006733,
  0.006085,   0.006085,    0.006085,    0.006085,
  0.005681,   0.005681,    0.005681,    0.005681,
  0.005445,   0.005445,    0.005445,    0.005445,
  0.005148,   0.005148,    0.005148,    0.005148,
  0.004982,   0.004982,    0.004982,    0.004982,
  0.005088,   0.005088,    0.005088,    0.005088,
  0.0051,     0.0051,      0.0051,      0.0051,
  0.004861,   0.004861,    0.004861,    0.004861,
  0.004854,   0.004854,    0.004854,    0.004854,
  0.004935,   0.004935,    0.004935,    0.004935,
  0.00486,    0.00486,     0.00486,     0.00486,
  0.004999,   0.004999,    0.004999,    0.004999,
  0.005163,   0.005163,    0.005163,    0.005163,
  0.004986,   0.004986,    0.004986,    0.004986,
  0.005012,   0.005012,    0.005012,    0.005012,
  0.005296,   0.005296,    0.005296,    0.005296,
  0.005465,   0.005465,    0.005465,    0.005465,
  0.005485,   0.005485,    0.005485,    0.005485,
  0.005636,   0.005636,    0.005636,    0.005636,
  0.006074,   0.006074,    0.006074,    0.006074,
  0.006522,   0.006522,    0.006522,    0.006522,
  0.00679,    0.00679,     0.00679,     0.00679,
  0.006956,   0.006956,    0.006956,    0.006956,
  0.007124,   0.007124,    0.007124,    0.007124,
  0.007544,   0.007544,    0.007544,    0.007544,
  0.008024,   0.008024,    0.008024,    0.008024,
  0.00821,    0.00821,     0.00821,     0.00821,
  0.008241,   0.008241,    0.008241,    0.008241,
  0.008238,   0.008238,    0.008238,    0.008238,
  0.008295,   0.008295,    0.008295,    0.008295,
  0.008388,   0.008388,    0.008388,    0.008388,
  0.008421,   0.008421,    0.008421,    0.008421,
  0.008423,   0.008423,    0.008423,    0.008423,
  0.008427,   0.008427,    0.008427,    0.008427,
  0.008397,   0.008397,    0.008397,    0.008397,
  0.008301,   0.008301,    0.008301,    0.008301,
  0.008205,   0.008205,    0.008205,    0.008205,
  0.008172,   0.008172,    0.008172,    0.008172,
  0.008305,   0.008305,    0.008305,    0.008305,
  0.008507,   0.008507,    0.008507,    0.008507,
  0.008572,   0.008572,    0.008572,    0.008572,
  0.008564,   0.008564,    0.008564,    0.008564,
  0.008526,   0.008526,    0.008526,    0.008526,
  0.008455,   0.008455,    0.008455,    0.008455,
  0.008299,   0.008299,    0.008299,    0.008299,
  0.008032,   0.008032,    0.008032,    0.008032,
  0.008006,   0.008006,    0.008006,    0.008006,
  0.007704,   0.007704,    0.007704,    0.007704,
  0.006603,   0.006603,    0.006603,    0.006603,
  0.005692,   0.005692,    0.005692,    0.005692,
  0.00517,    0.00517,     0.00517,     0.00517,
  0.004767,   0.004767,    0.004767,    0.004767,
  0.004584,   0.004584,    0.004584,    0.004584,
  0.004476,   0.004476,    0.004476,    0.004476,
  0.004437,   0.004437,    0.004437,    0.004437,
  0.004669,   0.004669,    0.004669,    0.004669,
  0.005559,   0.005559,    0.005559,    0.005559,
  0.006121,   0.006121,    0.006121,    0.006121,
  0.006164,   0.006164,    0.006164,    0.006164,
  0.006648,   0.006648,    0.006648,    0.006648,
  0.007522,   0.007522,    0.007522,    0.007522,
  0.007923,   0.007923,    0.007923,    0.007923,
  0.00786,    0.00786,     0.00786,     0.00786,
  0.007954,   0.007954,    0.007954,    0.007954,
  0.008436,   0.008436,    0.008436,    0.008436,
  0.008858,   0.008858,    0.008858,    0.008858,
  0.009047,   0.009047,    0.009047,    0.009047,
  0.009459,   0.009459,    0.009459,    0.009459,
  0.009881,   0.009881,    0.009881,    0.009881,
  0.01001,    0.01001,     0.01001,     0.01001,
  0.009897,   0.009897,    0.009897,    0.009897,
  0.009967,   0.009967,    0.009967,    0.009967,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.01022,    0.01022,     0.01022,     0.01022,
  0.01031,    0.01031,     0.01031,     0.01031,
  0.01035,    0.01035,     0.01035,     0.01035,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01024,    0.01024,     0.01024,     0.01024,
  0.01022,    0.01022,     0.01022,     0.01022,
  0.01014,    0.01014,     0.01014,     0.01014,
  0.01001,    0.01001,     0.01001,     0.01001,
  0.009865,   0.009865,    0.009865,    0.009865,
  0.009565,   0.009565,    0.009565,    0.009565,
  0.009295,   0.009295,    0.009295,    0.009295,
  0.009216,   0.009216,    0.009216,    0.009216,
  0.009137,   0.009137,    0.009137,    0.009137,
  0.009033,   0.009033,    0.009033,    0.009033,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.009138,   0.009138,    0.009138,    0.009138,
  0.009538,   0.009538,    0.009538,    0.009538,
  0.009979,   0.009979,    0.009979,    0.009979,
  0.01041,    0.01041,     0.01041,     0.01041,
  0.01079,    0.01079,     0.01079,     0.01079,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.00948,    0.00948,     0.00948,     0.00948,
  0.009003,   0.009003,    0.009003,    0.009003,
  0.008484,   0.008484,    0.008484,    0.008484,
  0.007951,   0.007951,    0.007951,    0.007951,
  0.007941,   0.007941,    0.007941,    0.007941,
  0.00847,    0.00847,     0.00847,     0.00847,
  0.008469,   0.008469,    0.008469,    0.008469,
  0.008253,   0.008253,    0.008253,    0.008253,
  0.008028,   0.008028,    0.008028,    0.008028,
  0.007983,   0.007983,    0.007983,    0.007983,
  0.007857,   0.007857,    0.007857,    0.007857,
  0.007628,   0.007628,    0.007628,    0.007628,
  0.007742,   0.007742,    0.007742,    0.007742,
  0.007872,   0.007872,    0.007872,    0.007872,
  0.007954,   0.007954,    0.007954,    0.007954,
  0.00834,    0.00834,     0.00834,     0.00834,
  0.008921,   0.008921,    0.008921,    0.008921,
  0.009234,   0.009234,    0.009234,    0.009234,
  0.009335,   0.009335,    0.009335,    0.009335,
  0.009333,   0.009333,    0.009333,    0.009333,
  0.009662,   0.009662,    0.009662,    0.009662,
  0.01013,    0.01013,     0.01013,     0.01013,
  0.01021,    0.01021,     0.01021,     0.01021,
  0.01012,    0.01012,     0.01012,     0.01012,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.01004,    0.01004,     0.01004,     0.01004,
  0.009955,   0.009955,    0.009955,    0.009955,
  0.009918,   0.009918,    0.009918,    0.009918,
  0.009971,   0.009971,    0.009971,    0.009971,
  0.009906,   0.009906,    0.009906,    0.009906,
  0.009856,   0.009856,    0.009856,    0.009856,
  0.009753,   0.009753,    0.009753,    0.009753,
  0.009577,   0.009577,    0.009577,    0.009577,
  0.009485,   0.009485,    0.009485,    0.009485,
  0.009481,   0.009481,    0.009481,    0.009481,
  0.0095,     0.0095,      0.0095,      0.0095,
  0.009366,   0.009366,    0.009366,    0.009366,
  0.009321,   0.009321,    0.009321,    0.009321,
  0.009396,   0.009396,    0.009396,    0.009396,
  0.009418,   0.009418,    0.009418,    0.009418,
  0.009477,   0.009477,    0.009477,    0.009477,
  0.009455,   0.009455,    0.009455,    0.009455,
  0.009509,   0.009509,    0.009509,    0.009509,
  0.009925,   0.009925,    0.009925,    0.009925,
  0.01041,    0.01041,     0.01041,     0.01041,
  0.01048,    0.01048,     0.01048,     0.01048,
  0.01012,    0.01012,     0.01012,     0.01012,
  0.009593,   0.009593,    0.009593,    0.009593,
  0.009115,   0.009115,    0.009115,    0.009115,
  0.008833,   0.008833,    0.008833,    0.008833,
  0.008799,   0.008799,    0.008799,    0.008799,
  0.009082,   0.009082,    0.009082,    0.009082,
  0.0091,     0.0091,      0.0091,      0.0091,
  0.008858,   0.008858,    0.008858,    0.008858,
  0.009098,   0.009098,    0.009098,    0.009098,
  0.009108,   0.009108,    0.009108,    0.009108,
  0.008812,   0.008812,    0.008812,    0.008812,
  0.008942,   0.008942,    0.008942,    0.008942,
  0.009002,   0.009002,    0.009002,    0.009002,
  0.008774,   0.008774,    0.008774,    0.008774,
  0.008711,   0.008711,    0.008711,    0.008711,
  0.008692,   0.008692,    0.008692,    0.008692,
  0.008536,   0.008536,    0.008536,    0.008536,
  0.008485,   0.008485,    0.008485,    0.008485,
  0.00885,    0.00885,     0.00885,     0.00885,
  0.009242,   0.009242,    0.009242,    0.009242,
  0.009103,   0.009103,    0.009103,    0.009103,
  0.008834,   0.008834,    0.008834,    0.008834,
  0.00862,    0.00862,     0.00862,     0.00862,
  0.008457,   0.008457,    0.008457,    0.008457,
  0.008493,   0.008493,    0.008493,    0.008493,
  0.008612,   0.008612,    0.008612,    0.008612,
  0.008756,   0.008756,    0.008756,    0.008756,
  0.008849,   0.008849,    0.008849,    0.008849,
  0.008903,   0.008903,    0.008903,    0.008903,
  0.008995,   0.008995,    0.008995,    0.008995,
  0.009015,   0.009015,    0.009015,    0.009015,
  0.008969,   0.008969,    0.008969,    0.008969,
  0.009011,   0.009011,    0.009011,    0.009011,
  0.009095,   0.009095,    0.009095,    0.009095,
  0.009132,   0.009132,    0.009132,    0.009132,
  0.009008,   0.009008,    0.009008,    0.009008,
  0.008779,   0.008779,    0.008779,    0.008779,
  0.008703,   0.008703,    0.008703,    0.008703,
  0.008654,   0.008654,    0.008654,    0.008654,
  0.00853,    0.00853,     0.00853,     0.00853,
  0.008432,   0.008432,    0.008432,    0.008432,
  0.008408,   0.008408,    0.008408,    0.008408,
  0.008384,   0.008384,    0.008384,    0.008384,
  0.008312,   0.008312,    0.008312,    0.008312,
  0.00836,    0.00836,     0.00836,     0.00836,
  0.00853,    0.00853,     0.00853,     0.00853,
  0.008754,   0.008754,    0.008754,    0.008754,
  0.009114,   0.009114,    0.009114,    0.009114,
  0.009565,   0.009565,    0.009565,    0.009565,
  0.009782,   0.009782,    0.009782,    0.009782,
  0.009576,   0.009576,    0.009576,    0.009576,
  0.009178,   0.009178,    0.009178,    0.009178,
  0.008989,   0.008989,    0.008989,    0.008989,
  0.008927,   0.008927,    0.008927,    0.008927,
  0.00877,    0.00877,     0.00877,     0.00877,
  0.008305,   0.008305,    0.008305,    0.008305,
  0.008366,   0.008366,    0.008366,    0.008366,
  0.008988,   0.008988,    0.008988,    0.008988,
  0.008865,   0.008865,    0.008865,    0.008865,
  0.008615,   0.008615,    0.008615,    0.008615,
  0.008585,   0.008585,    0.008585,    0.008585,
  0.008395,   0.008395,    0.008395,    0.008395,
  0.008162,   0.008162,    0.008162,    0.008162,
  0.008064,   0.008064,    0.008064,    0.008064,
  0.00852,    0.00852,     0.00852,     0.00852,
  0.009444,   0.009444,    0.009444,    0.009444,
  0.01005,    0.01005,     0.01005,     0.01005,
  0.01027,    0.01027,     0.01027,     0.01027,
  0.01054,    0.01054,     0.01054,     0.01054,
  0.01063,    0.01063,     0.01063,     0.01063,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.009523,   0.009523,    0.009523,    0.009523,
  0.009431,   0.009431,    0.009431,    0.009431,
  0.009372,   0.009372,    0.009372,    0.009372,
  0.00912,    0.00912,     0.00912,     0.00912,
  0.008936,   0.008936,    0.008936,    0.008936,
  0.00904,    0.00904,     0.00904,     0.00904,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.009019,   0.009019,    0.009019,    0.009019,
  0.008934,   0.008934,    0.008934,    0.008934,
  0.008828,   0.008828,    0.008828,    0.008828,
  0.008748,   0.008748,    0.008748,    0.008748,
  0.00876,    0.00876,     0.00876,     0.00876,
  0.008868,   0.008868,    0.008868,    0.008868,
  0.008945,   0.008945,    0.008945,    0.008945,
  0.009022,   0.009022,    0.009022,    0.009022,
  0.009032,   0.009032,    0.009032,    0.009032,
  0.009011,   0.009011,    0.009011,    0.009011,
  0.009033,   0.009033,    0.009033,    0.009033,
  0.009074,   0.009074,    0.009074,    0.009074,
  0.009121,   0.009121,    0.009121,    0.009121,
  0.009158,   0.009158,    0.009158,    0.009158,
  0.009268,   0.009268,    0.009268,    0.009268,
  0.009455,   0.009455,    0.009455,    0.009455,
  0.0097,     0.0097,      0.0097,      0.0097,
  0.01,       0.01,        0.01,        0.01,
  0.01022,    0.01022,     0.01022,     0.01022,
  0.01027,    0.01027,     0.01027,     0.01027,
  0.01033,    0.01033,     0.01033,     0.01033,
  0.0104,     0.0104,      0.0104,      0.0104,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01064,    0.01064,     0.01064,     0.01064,
  0.0106,     0.0106,      0.0106,      0.0106,
  0.01034,    0.01034,     0.01034,     0.01034,
  0.01034,    0.01034,     0.01034,     0.01034,
  0.01028,    0.01028,     0.01028,     0.01028,
  0.009946,   0.009946,    0.009946,    0.009946,
  0.009607,   0.009607,    0.009607,    0.009607,
  0.009418,   0.009418,    0.009418,    0.009418,
  0.009078,   0.009078,    0.009078,    0.009078,
  0.008598,   0.008598,    0.008598,    0.008598,
  0.008256,   0.008256,    0.008256,    0.008256,
  0.008118,   0.008118,    0.008118,    0.008118,
  0.00814,    0.00814,     0.00814,     0.00814,
  0.00819,    0.00819,     0.00819,     0.00819,
  0.008115,   0.008115,    0.008115,    0.008115,
  0.008076,   0.008076,    0.008076,    0.008076,
  0.007917,   0.007917,    0.007917,    0.007917,
  0.007917,   0.007917,    0.007917,    0.007917,
  0.008201,   0.008201,    0.008201,    0.008201,
  0.008332,   0.008332,    0.008332,    0.008332,
  0.008497,   0.008497,    0.008497,    0.008497,
  0.008694,   0.008694,    0.008694,    0.008694,
  0.008828,   0.008828,    0.008828,    0.008828,
  0.008929,   0.008929,    0.008929,    0.008929,
  0.009002,   0.009002,    0.009002,    0.009002,
  0.009108,   0.009108,    0.009108,    0.009108,
  0.00918,    0.00918,     0.00918,     0.00918,
  0.009218,   0.009218,    0.009218,    0.009218,
  0.009284,   0.009284,    0.009284,    0.009284,
  0.009322,   0.009322,    0.009322,    0.009322,
  0.009329,   0.009329,    0.009329,    0.009329,
  0.009337,   0.009337,    0.009337,    0.009337,
  0.009372,   0.009372,    0.009372,    0.009372,
  0.009408,   0.009408,    0.009408,    0.009408,
  0.009415,   0.009415,    0.009415,    0.009415,
  0.009455,   0.009455,    0.009455,    0.009455,
  0.009487,   0.009487,    0.009487,    0.009487,
  0.009487,   0.009487,    0.009487,    0.009487,
  0.009546,   0.009546,    0.009546,    0.009546,
  0.009652,   0.009652,    0.009652,    0.009652,
  0.009751,   0.009751,    0.009751,    0.009751,
  0.009788,   0.009788,    0.009788,    0.009788,
  0.009678,   0.009678,    0.009678,    0.009678,
  0.009446,   0.009446,    0.009446,    0.009446,
  0.009149,   0.009149,    0.009149,    0.009149,
  0.00883,    0.00883,     0.00883,     0.00883,
  0.008546,   0.008546,    0.008546,    0.008546,
  0.008293,   0.008293,    0.008293,    0.008293,
  0.008043,   0.008043,    0.008043,    0.008043,
  0.008043,   0.008043,    0.008043,    0.008043,
  0.00814,    0.00814,     0.00814,     0.00814,
  0.008087,   0.008087,    0.008087,    0.008087,
  0.007873,   0.007873,    0.007873,    0.007873,
  0.007712,   0.007712,    0.007712,    0.007712,
  0.007744,   0.007744,    0.007744,    0.007744,
  0.007717,   0.007717,    0.007717,    0.007717,
  0.005882,   0.005882,    0.005882,    0.005882,
  0.005586,   0.005586,    0.005586,    0.005586,
  0.006817,   0.006817,    0.006817,    0.006817,
  0.006447,   0.006447,    0.006447,    0.006447,
  0.00625,    0.00625,     0.00625,     0.00625,
  0.006014,   0.006014,    0.006014,    0.006014,
  0.005815,   0.005815,    0.005815,    0.005815,
  0.005815,   0.005815,    0.005815,    0.005815,
  0.005694,   0.005694,    0.005694,    0.005694,
  0.005941,   0.005941,    0.005941,    0.005941,
  0.006534,   0.006534,    0.006534,    0.006534,
  0.006791,   0.006791,    0.006791,    0.006791,
  0.007032,   0.007032,    0.007032,    0.007032,
  0.007221,   0.007221,    0.007221,    0.007221,
  0.007318,   0.007318,    0.007318,    0.007318,
  0.00728,    0.00728,     0.00728,     0.00728,
  0.007319,   0.007319,    0.007319,    0.007319,
  0.00754,    0.00754,     0.00754,     0.00754,
  0.007697,   0.007697,    0.007697,    0.007697,
  0.007925,   0.007925,    0.007925,    0.007925,
  0.00812,    0.00812,     0.00812,     0.00812,
  0.008183,   0.008183,    0.008183,    0.008183,
  0.008191,   0.008191,    0.008191,    0.008191,
  0.008198,   0.008198,    0.008198,    0.008198,
  0.008205,   0.008205,    0.008205,    0.008205,
  0.008156,   0.008156,    0.008156,    0.008156,
  0.008108,   0.008108,    0.008108,    0.008108,
  0.008084,   0.008084,    0.008084,    0.008084,
  0.008115,   0.008115,    0.008115,    0.008115,
  0.008186,   0.008186,    0.008186,    0.008186,
  0.008225,   0.008225,    0.008225,    0.008225,
  0.008266,   0.008266,    0.008266,    0.008266,
  0.008373,   0.008373,    0.008373,    0.008373,
  0.008528,   0.008528,    0.008528,    0.008528,
  0.008624,   0.008624,    0.008624,    0.008624,
  0.008496,   0.008496,    0.008496,    0.008496,
  0.00825,    0.00825,     0.00825,     0.00825,
  0.008096,   0.008096,    0.008096,    0.008096,
  0.00816,    0.00816,     0.00816,     0.00816,
  0.008404,   0.008404,    0.008404,    0.008404,
  0.008616,   0.008616,    0.008616,    0.008616,
  0.008654,   0.008654,    0.008654,    0.008654,
  0.008832,   0.008832,    0.008832,    0.008832,
  0.009147,   0.009147,    0.009147,    0.009147,
  0.00896,    0.00896,     0.00896,     0.00896,
  0.008234,   0.008234,    0.008234,    0.008234,
  0.007728,   0.007728,    0.007728,    0.007728,
  0.007601,   0.007601,    0.007601,    0.007601,
  0.006719,   0.006719,    0.006719,    0.006719,
  0.006659,   0.006659,    0.006659,    0.006659,
  0.007131,   0.007131,    0.007131,    0.007131,
  0.006907,   0.006907,    0.006907,    0.006907,
  0.007003,   0.007003,    0.007003,    0.007003,
  0.007038,   0.007038,    0.007038,    0.007038,
  0.007075,   0.007075,    0.007075,    0.007075,
  0.007234,   0.007234,    0.007234,    0.007234,
  0.00705,    0.00705,     0.00705,     0.00705,
  0.007033,   0.007033,    0.007033,    0.007033,
  0.007512,   0.007512,    0.007512,    0.007512,
  0.007854,   0.007854,    0.007854,    0.007854,
  0.008229,   0.008229,    0.008229,    0.008229,
  0.008547,   0.008547,    0.008547,    0.008547,
  0.008711,   0.008711,    0.008711,    0.008711,
  0.008813,   0.008813,    0.008813,    0.008813,
  0.008888,   0.008888,    0.008888,    0.008888,
  0.008882,   0.008882,    0.008882,    0.008882,
  0.008763,   0.008763,    0.008763,    0.008763,
  0.008825,   0.008825,    0.008825,    0.008825,
  0.008965,   0.008965,    0.008965,    0.008965,
  0.008975,   0.008975,    0.008975,    0.008975,
  0.008953,   0.008953,    0.008953,    0.008953,
  0.008958,   0.008958,    0.008958,    0.008958,
  0.008964,   0.008964,    0.008964,    0.008964,
  0.008885,   0.008885,    0.008885,    0.008885,
  0.008833,   0.008833,    0.008833,    0.008833,
  0.008807,   0.008807,    0.008807,    0.008807,
  0.008787,   0.008787,    0.008787,    0.008787,
  0.00883,    0.00883,     0.00883,     0.00883,
  0.008868,   0.008868,    0.008868,    0.008868,
  0.008887,   0.008887,    0.008887,    0.008887,
  0.009086,   0.009086,    0.009086,    0.009086,
  0.009394,   0.009394,    0.009394,    0.009394,
  0.009568,   0.009568,    0.009568,    0.009568,
  0.00957,    0.00957,     0.00957,     0.00957,
  0.009666,   0.009666,    0.009666,    0.009666,
  0.009965,   0.009965,    0.009965,    0.009965,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01062,    0.01062,     0.01062,     0.01062,
  0.01088,    0.01088,     0.01088,     0.01088,
  0.01095,    0.01095,     0.01095,     0.01095,
  0.0108,     0.0108,      0.0108,      0.0108,
  0.01078,    0.01078,     0.01078,     0.01078,
  0.0105,     0.0105,      0.0105,      0.0105,
  0.008655,   0.008655,    0.008655,    0.008655,
  0.007155,   0.007155,    0.007155,    0.007155,
  0.007612,   0.007612,    0.007612,    0.007612,
  0.007504,   0.007504,    0.007504,    0.007504,
  0.007766,   0.007766,    0.007766,    0.007766,
  0.0085,     0.0085,      0.0085,      0.0085,
  0.008679,   0.008679,    0.008679,    0.008679,
  0.009085,   0.009085,    0.009085,    0.009085,
  0.00941,    0.00941,     0.00941,     0.00941,
  0.009491,   0.009491,    0.009491,    0.009491,
  0.0095,     0.0095,      0.0095,      0.0095,
  0.009264,   0.009264,    0.009264,    0.009264,
  0.009136,   0.009136,    0.009136,    0.009136,
  0.009463,   0.009463,    0.009463,    0.009463,
  0.009447,   0.009447,    0.009447,    0.009447,
  0.008677,   0.008677,    0.008677,    0.008677,
  0.007922,   0.007922,    0.007922,    0.007922,
  0.007791,   0.007791,    0.007791,    0.007791,
  0.007793,   0.007793,    0.007793,    0.007793,
  0.007826,   0.007826,    0.007826,    0.007826,
  0.007917,   0.007917,    0.007917,    0.007917,
  0.0081,     0.0081,      0.0081,      0.0081,
  0.008326,   0.008326,    0.008326,    0.008326,
  0.008496,   0.008496,    0.008496,    0.008496,
  0.008559,   0.008559,    0.008559,    0.008559,
  0.008565,   0.008565,    0.008565,    0.008565,
  0.008546,   0.008546,    0.008546,    0.008546,
  0.008526,   0.008526,    0.008526,    0.008526,
  0.008476,   0.008476,    0.008476,    0.008476,
  0.008401,   0.008401,    0.008401,    0.008401,
  0.008327,   0.008327,    0.008327,    0.008327,
  0.008285,   0.008285,    0.008285,    0.008285,
  0.008331,   0.008331,    0.008331,    0.008331,
  0.008394,   0.008394,    0.008394,    0.008394,
  0.008485,   0.008485,    0.008485,    0.008485,
  0.008673,   0.008673,    0.008673,    0.008673,
  0.008913,   0.008913,    0.008913,    0.008913,
  0.0091,     0.0091,      0.0091,      0.0091,
  0.009317,   0.009317,    0.009317,    0.009317,
  0.009455,   0.009455,    0.009455,    0.009455,
  0.009624,   0.009624,    0.009624,    0.009624,
  0.01016,    0.01016,     0.01016,     0.01016,
  0.01065,    0.01065,     0.01065,     0.01065,
  0.01081,    0.01081,     0.01081,     0.01081,
  0.01063,    0.01063,     0.01063,     0.01063,
  0.01063,    0.01063,     0.01063,     0.01063,
  0.01075,    0.01075,     0.01075,     0.01075,
  0.009271,   0.009271,    0.009271,    0.009271,
  0.007826,   0.007826,    0.007826,    0.007826,
  0.007485,   0.007485,    0.007485,    0.007485,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.006601,   0.006601,    0.006601,    0.006601,
  0.00702,    0.00702,     0.00702,     0.00702,
  0.007304,   0.007304,    0.007304,    0.007304,
  0.006846,   0.006846,    0.006846,    0.006846,
  0.007222,   0.007222,    0.007222,    0.007222,
  0.007318,   0.007318,    0.007318,    0.007318,
  0.007603,   0.007603,    0.007603,    0.007603,
  0.008305,   0.008305,    0.008305,    0.008305,
  0.008341,   0.008341,    0.008341,    0.008341,
  0.008528,   0.008528,    0.008528,    0.008528,
  0.009128,   0.009128,    0.009128,    0.009128,
  0.009215,   0.009215,    0.009215,    0.009215,
  0.009146,   0.009146,    0.009146,    0.009146,
  0.008967,   0.008967,    0.008967,    0.008967,
  0.008828,   0.008828,    0.008828,    0.008828,
  0.008756,   0.008756,    0.008756,    0.008756,
  0.008689,   0.008689,    0.008689,    0.008689,
  0.008715,   0.008715,    0.008715,    0.008715,
  0.008817,   0.008817,    0.008817,    0.008817,
  0.009096,   0.009096,    0.009096,    0.009096,
  0.009345,   0.009345,    0.009345,    0.009345,
  0.009435,   0.009435,    0.009435,    0.009435,
  0.009412,   0.009412,    0.009412,    0.009412,
  0.009388,   0.009388,    0.009388,    0.009388,
  0.009475,   0.009475,    0.009475,    0.009475,
  0.009641,   0.009641,    0.009641,    0.009641,
  0.009753,   0.009753,    0.009753,    0.009753,
  0.009725,   0.009725,    0.009725,    0.009725,
  0.009757,   0.009757,    0.009757,    0.009757,
  0.009936,   0.009936,    0.009936,    0.009936,
  0.01008,    0.01008,     0.01008,     0.01008,
  0.01026,    0.01026,     0.01026,     0.01026,
  0.01043,    0.01043,     0.01043,     0.01043,
  0.01048,    0.01048,     0.01048,     0.01048,
  0.01051,    0.01051,     0.01051,     0.01051,
  0.0106,     0.0106,      0.0106,      0.0106,
  0.01076,    0.01076,     0.01076,     0.01076,
  0.01088,    0.01088,     0.01088,     0.01088,
  0.01085,    0.01085,     0.01085,     0.01085,
  0.0111,     0.0111,      0.0111,      0.0111,
  0.01137,    0.01137,     0.01137,     0.01137,
  0.01106,    0.01106,     0.01106,     0.01106,
  0.01077,    0.01077,     0.01077,     0.01077,
  0.01071,    0.01071,     0.01071,     0.01071,
  0.01058,    0.01058,     0.01058,     0.01058,
  0.01038,    0.01038,     0.01038,     0.01038,
  0.009907,   0.009907,    0.009907,    0.009907,
  0.00915,    0.00915,     0.00915,     0.00915,
  0.006818,   0.006818,    0.006818,    0.006818,
  0.005489,   0.005489,    0.005489,    0.005489,
  0.006237,   0.006237,    0.006237,    0.006237,
  0.006267,   0.006267,    0.006267,    0.006267,
  0.006335,   0.006335,    0.006335,    0.006335,
  0.006617,   0.006617,    0.006617,    0.006617,
  0.006835,   0.006835,    0.006835,    0.006835,
  0.007024,   0.007024,    0.007024,    0.007024,
  0.006871,   0.006871,    0.006871,    0.006871,
  0.007003,   0.007003,    0.007003,    0.007003,
  0.007541,   0.007541,    0.007541,    0.007541,
  0.007824,   0.007824,    0.007824,    0.007824,
  0.0082,     0.0082,      0.0082,      0.0082,
  0.008605,   0.008605,    0.008605,    0.008605,
  0.008916,   0.008916,    0.008916,    0.008916,
  0.009165,   0.009165,    0.009165,    0.009165,
  0.009383,   0.009383,    0.009383,    0.009383,
  0.009604,   0.009604,    0.009604,    0.009604,
  0.009761,   0.009761,    0.009761,    0.009761,
  0.01001,    0.01001,     0.01001,     0.01001,
  0.01026,    0.01026,     0.01026,     0.01026,
  0.01036,    0.01036,     0.01036,     0.01036,
  0.01036,    0.01036,     0.01036,     0.01036,
  0.01036,    0.01036,     0.01036,     0.01036,
  0.01033,    0.01033,     0.01033,     0.01033,
  0.01018,    0.01018,     0.01018,     0.01018,
  0.01001,    0.01001,     0.01001,     0.01001,
  0.009867,   0.009867,    0.009867,    0.009867,
  0.009785,   0.009785,    0.009785,    0.009785,
  0.009767,   0.009767,    0.009767,    0.009767,
  0.00983,    0.00983,     0.00983,     0.00983,
  0.009854,   0.009854,    0.009854,    0.009854,
  0.009848,   0.009848,    0.009848,    0.009848,
  0.009838,   0.009838,    0.009838,    0.009838,
  0.009824,   0.009824,    0.009824,    0.009824,
  0.009714,   0.009714,    0.009714,    0.009714,
  0.009484,   0.009484,    0.009484,    0.009484,
  0.009408,   0.009408,    0.009408,    0.009408,
  0.009556,   0.009556,    0.009556,    0.009556,
  0.009648,   0.009648,    0.009648,    0.009648,
  0.009616,   0.009616,    0.009616,    0.009616,
  0.009657,   0.009657,    0.009657,    0.009657,
  0.009935,   0.009935,    0.009935,    0.009935,
  0.01029,    0.01029,     0.01029,     0.01029,
  0.01029,    0.01029,     0.01029,     0.01029,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.009796,   0.009796,    0.009796,    0.009796,
  0.009289,   0.009289,    0.009289,    0.009289,
  0.007972,   0.007972,    0.007972,    0.007972,
  0.007801,   0.007801,    0.007801,    0.007801,
  0.008821,   0.008821,    0.008821,    0.008821,
  0.008821,   0.008821,    0.008821,    0.008821,
  0.008906,   0.008906,    0.008906,    0.008906,
  0.009447,   0.009447,    0.009447,    0.009447,
  0.009564,   0.009564,    0.009564,    0.009564,
  0.009429,   0.009429,    0.009429,    0.009429,
  0.009054,   0.009054,    0.009054,    0.009054,
  0.008964,   0.008964,    0.008964,    0.008964,
  0.009295,   0.009295,    0.009295,    0.009295,
  0.009216,   0.009216,    0.009216,    0.009216,
  0.009114,   0.009114,    0.009114,    0.009114,
  0.009178,   0.009178,    0.009178,    0.009178,
  0.009157,   0.009157,    0.009157,    0.009157,
  0.00896,    0.00896,     0.00896,     0.00896,
  0.008859,   0.008859,    0.008859,    0.008859,
  0.008854,   0.008854,    0.008854,    0.008854,
  0.008817,   0.008817,    0.008817,    0.008817,
  0.008987,   0.008987,    0.008987,    0.008987,
  0.009153,   0.009153,    0.009153,    0.009153,
  0.009081,   0.009081,    0.009081,    0.009081,
  0.008875,   0.008875,    0.008875,    0.008875,
  0.008597,   0.008597,    0.008597,    0.008597,
  0.008552,   0.008552,    0.008552,    0.008552,
  0.008704,   0.008704,    0.008704,    0.008704,
  0.008807,   0.008807,    0.008807,    0.008807,
  0.008885,   0.008885,    0.008885,    0.008885,
  0.008995,   0.008995,    0.008995,    0.008995,
  0.009116,   0.009116,    0.009116,    0.009116,
  0.009075,   0.009075,    0.009075,    0.009075,
  0.008939,   0.008939,    0.008939,    0.008939,
  0.00898,    0.00898,     0.00898,     0.00898,
  0.00915,    0.00915,     0.00915,     0.00915,
  0.00946,    0.00946,     0.00946,     0.00946,
  0.009776,   0.009776,    0.009776,    0.009776,
  0.009814,   0.009814,    0.009814,    0.009814,
  0.009744,   0.009744,    0.009744,    0.009744,
  0.009805,   0.009805,    0.009805,    0.009805,
  0.009997,   0.009997,    0.009997,    0.009997,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.01028,    0.01028,     0.01028,     0.01028,
  0.01057,    0.01057,     0.01057,     0.01057,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.01034,    0.01034,     0.01034,     0.01034,
  0.01016,    0.01016,     0.01016,     0.01016,
  0.01027,    0.01027,     0.01027,     0.01027,
  0.009461,   0.009461,    0.009461,    0.009461,
  0.009268,   0.009268,    0.009268,    0.009268,
  0.01013,    0.01013,     0.01013,     0.01013,
  0.01021,    0.01021,     0.01021,     0.01021,
  0.01048,    0.01048,     0.01048,     0.01048,
  0.01078,    0.01078,     0.01078,     0.01078,
  0.01085,    0.01085,     0.01085,     0.01085,
  0.01096,    0.01096,     0.01096,     0.01096,
  0.01078,    0.01078,     0.01078,     0.01078,
  0.01081,    0.01081,     0.01081,     0.01081,
  0.01093,    0.01093,     0.01093,     0.01093,
  0.01066,    0.01066,     0.01066,     0.01066,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01027,    0.01027,     0.01027,     0.01027,
  0.009938,   0.009938,    0.009938,    0.009938,
  0.009528,   0.009528,    0.009528,    0.009528,
  0.009325,   0.009325,    0.009325,    0.009325,
  0.009195,   0.009195,    0.009195,    0.009195,
  0.009266,   0.009266,    0.009266,    0.009266,
  0.009546,   0.009546,    0.009546,    0.009546,
  0.009404,   0.009404,    0.009404,    0.009404,
  0.009162,   0.009162,    0.009162,    0.009162,
  0.00914,    0.00914,     0.00914,     0.00914,
  0.009225,   0.009225,    0.009225,    0.009225,
  0.009284,   0.009284,    0.009284,    0.009284,
  0.009096,   0.009096,    0.009096,    0.009096,
  0.008809,   0.008809,    0.008809,    0.008809,
  0.008502,   0.008502,    0.008502,    0.008502,
  0.008383,   0.008383,    0.008383,    0.008383,
  0.008478,   0.008478,    0.008478,    0.008478,
  0.00859,    0.00859,     0.00859,     0.00859,
  0.008684,   0.008684,    0.008684,    0.008684,
  0.009036,   0.009036,    0.009036,    0.009036,
  0.009735,   0.009735,    0.009735,    0.009735,
  0.01051,    0.01051,     0.01051,     0.01051,
  0.01091,    0.01091,     0.01091,     0.01091,
  0.01092,    0.01092,     0.01092,     0.01092,
  0.01091,    0.01091,     0.01091,     0.01091,
  0.01106,    0.01106,     0.01106,     0.01106,
  0.01131,    0.01131,     0.01131,     0.01131,
  0.01144,    0.01144,     0.01144,     0.01144,
  0.01135,    0.01135,     0.01135,     0.01135,
  0.01124,    0.01124,     0.01124,     0.01124,
  0.01118,    0.01118,     0.01118,     0.01118,
  0.01072,    0.01072,     0.01072,     0.01072,
  0.009471,   0.009471,    0.009471,    0.009471,
  0.008142,   0.008142,    0.008142,    0.008142,
  0.007417,   0.007417,    0.007417,    0.007417,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006184,   0.006184,    0.006184,    0.006184,
  0.006939,   0.006939,    0.006939,    0.006939,
  0.007258,   0.007258,    0.007258,    0.007258,
  0.007839,   0.007839,    0.007839,    0.007839,
  0.0086,     0.0086,      0.0086,      0.0086,
  0.009169,   0.009169,    0.009169,    0.009169,
  0.009358,   0.009358,    0.009358,    0.009358,
  0.009123,   0.009123,    0.009123,    0.009123,
  0.00917,    0.00917,     0.00917,     0.00917,
  0.009531,   0.009531,    0.009531,    0.009531,
  0.009612,   0.009612,    0.009612,    0.009612,
  0.009791,   0.009791,    0.009791,    0.009791,
  0.01001,    0.01001,     0.01001,     0.01001,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.009932,   0.009932,    0.009932,    0.009932,
  0.009839,   0.009839,    0.009839,    0.009839,
  0.009638,   0.009638,    0.009638,    0.009638,
  0.009323,   0.009323,    0.009323,    0.009323,
  0.009432,   0.009432,    0.009432,    0.009432,
  0.009485,   0.009485,    0.009485,    0.009485,
  0.009435,   0.009435,    0.009435,    0.009435,
  0.009439,   0.009439,    0.009439,    0.009439,
  0.009388,   0.009388,    0.009388,    0.009388,
  0.009475,   0.009475,    0.009475,    0.009475,
  0.00953,    0.00953,     0.00953,     0.00953,
  0.009613,   0.009613,    0.009613,    0.009613,
  0.009669,   0.009669,    0.009669,    0.009669,
  0.009644,   0.009644,    0.009644,    0.009644,
  0.009628,   0.009628,    0.009628,    0.009628,
  0.009473,   0.009473,    0.009473,    0.009473,
  0.009253,   0.009253,    0.009253,    0.009253,
  0.009111,   0.009111,    0.009111,    0.009111,
  0.008937,   0.008937,    0.008937,    0.008937,
  0.00878,    0.00878,     0.00878,     0.00878,
  0.008655,   0.008655,    0.008655,    0.008655,
  0.008437,   0.008437,    0.008437,    0.008437,
  0.008096,   0.008096,    0.008096,    0.008096,
  0.007916,   0.007916,    0.007916,    0.007916,
  0.008043,   0.008043,    0.008043,    0.008043,
  0.008215,   0.008215,    0.008215,    0.008215,
  0.008389,   0.008389,    0.008389,    0.008389,
  0.008583,   0.008583,    0.008583,    0.008583,
  0.008398,   0.008398,    0.008398,    0.008398,
  0.008053,   0.008053,    0.008053,    0.008053,
  0.007795,   0.007795,    0.007795,    0.007795,
  0.00699,    0.00699,     0.00699,     0.00699,
  0.006711,   0.006711,    0.006711,    0.006711,
  0.006255,   0.006255,    0.006255,    0.006255,
  0.006122,   0.006122,    0.006122,    0.006122,
  0.00669,    0.00669,     0.00669,     0.00669,
  0.006447,   0.006447,    0.006447,    0.006447,
  0.006307,   0.006307,    0.006307,    0.006307,
  0.006296,   0.006296,    0.006296,    0.006296,
  0.006399,   0.006399,    0.006399,    0.006399,
  0.006761,   0.006761,    0.006761,    0.006761,
  0.006812,   0.006812,    0.006812,    0.006812,
  0.007003,   0.007003,    0.007003,    0.007003,
  0.007512,   0.007512,    0.007512,    0.007512,
  0.007651,   0.007651,    0.007651,    0.007651,
  0.007825,   0.007825,    0.007825,    0.007825,
  0.007976,   0.007976,    0.007976,    0.007976,
  0.007952,   0.007952,    0.007952,    0.007952,
  0.007899,   0.007899,    0.007899,    0.007899,
  0.007878,   0.007878,    0.007878,    0.007878,
  0.007968,   0.007968,    0.007968,    0.007968,
  0.008074,   0.008074,    0.008074,    0.008074,
  0.008352,   0.008352,    0.008352,    0.008352,
  0.00865,    0.00865,     0.00865,     0.00865,
  0.008843,   0.008843,    0.008843,    0.008843,
  0.009033,   0.009033,    0.009033,    0.009033,
  0.009144,   0.009144,    0.009144,    0.009144,
  0.009229,   0.009229,    0.009229,    0.009229,
  0.009283,   0.009283,    0.009283,    0.009283,
  0.009338,   0.009338,    0.009338,    0.009338,
  0.009365,   0.009365,    0.009365,    0.009365,
  0.009396,   0.009396,    0.009396,    0.009396,
  0.009464,   0.009464,    0.009464,    0.009464,
  0.009499,   0.009499,    0.009499,    0.009499,
  0.00955,    0.00955,     0.00955,     0.00955,
  0.009652,   0.009652,    0.009652,    0.009652,
  0.009725,   0.009725,    0.009725,    0.009725,
  0.009709,   0.009709,    0.009709,    0.009709,
  0.009687,   0.009687,    0.009687,    0.009687,
  0.009633,   0.009633,    0.009633,    0.009633,
  0.009529,   0.009529,    0.009529,    0.009529,
  0.009713,   0.009713,    0.009713,    0.009713,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.0102,     0.0102,      0.0102,      0.0102,
  0.01012,    0.01012,     0.01012,     0.01012,
  0.01007,    0.01007,     0.01007,     0.01007,
  0.01022,    0.01022,     0.01022,     0.01022,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.009934,   0.009934,    0.009934,    0.009934,
  0.0089,     0.0089,      0.0089,      0.0089,
  0.008738,   0.008738,    0.008738,    0.008738,
  0.009405,   0.009405,    0.009405,    0.009405,
  0.009442,   0.009442,    0.009442,    0.009442,
  0.009452,   0.009452,    0.009452,    0.009452,
  0.009519,   0.009519,    0.009519,    0.009519,
  0.009599,   0.009599,    0.009599,    0.009599,
  0.009536,   0.009536,    0.009536,    0.009536,
  0.009054,   0.009054,    0.009054,    0.009054,
  0.009032,   0.009032,    0.009032,    0.009032,
  0.009396,   0.009396,    0.009396,    0.009396,
  0.009346,   0.009346,    0.009346,    0.009346,
  0.009496,   0.009496,    0.009496,    0.009496,
  0.00965,    0.00965,     0.00965,     0.00965,
  0.009679,   0.009679,    0.009679,    0.009679,
  0.00953,    0.00953,     0.00953,     0.00953,
  0.009208,   0.009208,    0.009208,    0.009208,
  0.009223,   0.009223,    0.009223,    0.009223,
  0.009467,   0.009467,    0.009467,    0.009467,
  0.009866,   0.009866,    0.009866,    0.009866,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.01045,    0.01045,     0.01045,     0.01045,
  0.0106,     0.0106,      0.0106,      0.0106,
  0.01078,    0.01078,     0.01078,     0.01078,
  0.01097,    0.01097,     0.01097,     0.01097,
  0.01094,    0.01094,     0.01094,     0.01094,
  0.01079,    0.01079,     0.01079,     0.01079,
  0.01069,    0.01069,     0.01069,     0.01069,
  0.01069,    0.01069,     0.01069,     0.01069,
  0.01079,    0.01079,     0.01079,     0.01079,
  0.01073,    0.01073,     0.01073,     0.01073,
  0.01049,    0.01049,     0.01049,     0.01049,
  0.01037,    0.01037,     0.01037,     0.01037,
  0.01027,    0.01027,     0.01027,     0.01027,
  0.01017,    0.01017,     0.01017,     0.01017,
  0.0101,     0.0101,      0.0101,      0.0101,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.009963,   0.009963,    0.009963,    0.009963,
  0.009713,   0.009713,    0.009713,    0.009713,
  0.00922,    0.00922,     0.00922,     0.00922,
  0.00897,    0.00897,     0.00897,     0.00897,
  0.008743,   0.008743,    0.008743,    0.008743,
  0.008552,   0.008552,    0.008552,    0.008552,
  0.008611,   0.008611,    0.008611,    0.008611,
  0.008265,   0.008265,    0.008265,    0.008265,
  0.007795,   0.007795,    0.007795,    0.007795,
  0.007574,   0.007574,    0.007574,    0.007574,
  0.007205,   0.007205,    0.007205,    0.007205,
  0.005983,   0.005983,    0.005983,    0.005983,
  0.005848,   0.005848,    0.005848,    0.005848,
  0.006721,   0.006721,    0.006721,    0.006721,
  0.006629,   0.006629,    0.006629,    0.006629,
  0.006664,   0.006664,    0.006664,    0.006664,
  0.006977,   0.006977,    0.006977,    0.006977,
  0.007227,   0.007227,    0.007227,    0.007227,
  0.007447,   0.007447,    0.007447,    0.007447,
  0.007291,   0.007291,    0.007291,    0.007291,
  0.00736,    0.00736,     0.00736,     0.00736,
  0.007659,   0.007659,    0.007659,    0.007659,
  0.007538,   0.007538,    0.007538,    0.007538,
  0.007464,   0.007464,    0.007464,    0.007464,
  0.007485,   0.007485,    0.007485,    0.007485,
  0.0075,     0.0075,      0.0075,      0.0075,
  0.007457,   0.007457,    0.007457,    0.007457,
  0.007444,   0.007444,    0.007444,    0.007444,
  0.00754,    0.00754,     0.00754,     0.00754,
  0.007503,   0.007503,    0.007503,    0.007503,
  0.007586,   0.007586,    0.007586,    0.007586,
  0.007689,   0.007689,    0.007689,    0.007689,
  0.007705,   0.007705,    0.007705,    0.007705,
  0.007807,   0.007807,    0.007807,    0.007807,
  0.007745,   0.007745,    0.007745,    0.007745,
  0.007481,   0.007481,    0.007481,    0.007481,
  0.007213,   0.007213,    0.007213,    0.007213,
  0.006998,   0.006998,    0.006998,    0.006998,
  0.00685,    0.00685,     0.00685,     0.00685,
  0.006881,   0.006881,    0.006881,    0.006881,
  0.007039,   0.007039,    0.007039,    0.007039,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007113,   0.007113,    0.007113,    0.007113,
  0.007288,   0.007288,    0.007288,    0.007288,
  0.007761,   0.007761,    0.007761,    0.007761,
  0.008351,   0.008351,    0.008351,    0.008351,
  0.00905,    0.00905,     0.00905,     0.00905,
  0.009607,   0.009607,    0.009607,    0.009607,
  0.009902,   0.009902,    0.009902,    0.009902,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.01059,    0.01059,     0.01059,     0.01059,
  0.01081,    0.01081,     0.01081,     0.01081,
  0.01092,    0.01092,     0.01092,     0.01092,
  0.01106,    0.01106,     0.01106,     0.01106,
  0.01118,    0.01118,     0.01118,     0.01118,
  0.01098,    0.01098,     0.01098,     0.01098,
  0.01068,    0.01068,     0.01068,     0.01068,
  0.01049,    0.01049,     0.01049,     0.01049,
  0.01042,    0.01042,     0.01042,     0.01042,
  0.009198,   0.009198,    0.009198,    0.009198,
  0.008553,   0.008553,    0.008553,    0.008553,
  0.009332,   0.009332,    0.009332,    0.009332,
  0.009368,   0.009368,    0.009368,    0.009368,
  0.009451,   0.009451,    0.009451,    0.009451,
  0.009852,   0.009852,    0.009852,    0.009852,
  0.01004,    0.01004,     0.01004,     0.01004,
  0.009935,   0.009935,    0.009935,    0.009935,
  0.009442,   0.009442,    0.009442,    0.009442,
  0.009241,   0.009241,    0.009241,    0.009241,
  0.009264,   0.009264,    0.009264,    0.009264,
  0.00899,    0.00899,     0.00899,     0.00899,
  0.008894,   0.008894,    0.008894,    0.008894,
  0.008904,   0.008904,    0.008904,    0.008904,
  0.008887,   0.008887,    0.008887,    0.008887,
  0.008757,   0.008757,    0.008757,    0.008757,
  0.008633,   0.008633,    0.008633,    0.008633,
  0.00866,    0.00866,     0.00866,     0.00866,
  0.008627,   0.008627,    0.008627,    0.008627,
  0.008639,   0.008639,    0.008639,    0.008639,
  0.008754,   0.008754,    0.008754,    0.008754,
  0.008513,   0.008513,    0.008513,    0.008513,
  0.00807,    0.00807,     0.00807,     0.00807,
  0.008053,   0.008053,    0.008053,    0.008053,
  0.00818,    0.00818,     0.00818,     0.00818,
  0.008156,   0.008156,    0.008156,    0.008156,
  0.008084,   0.008084,    0.008084,    0.008084,
  0.007871,   0.007871,    0.007871,    0.007871,
  0.007535,   0.007535,    0.007535,    0.007535,
  0.007405,   0.007405,    0.007405,    0.007405,
  0.007512,   0.007512,    0.007512,    0.007512,
  0.007682,   0.007682,    0.007682,    0.007682,
  0.008088,   0.008088,    0.008088,    0.008088,
  0.008658,   0.008658,    0.008658,    0.008658,
  0.009242,   0.009242,    0.009242,    0.009242,
  0.00975,    0.00975,     0.00975,     0.00975,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01068,    0.01068,     0.01068,     0.01068,
  0.01106,    0.01106,     0.01106,     0.01106,
  0.01126,    0.01126,     0.01126,     0.01126,
  0.01102,    0.01102,     0.01102,     0.01102,
  0.01095,    0.01095,     0.01095,     0.01095,
  0.0113,     0.0113,      0.0113,      0.0113,
  0.01124,    0.01124,     0.01124,     0.01124,
  0.0111,     0.0111,      0.0111,      0.0111,
  0.01107,    0.01107,     0.01107,     0.01107,
  0.01104,    0.01104,     0.01104,     0.01104,
  0.0102,     0.0102,      0.0102,      0.0102,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.01081,    0.01081,     0.01081,     0.01081,
  0.01081,    0.01081,     0.01081,     0.01081,
  0.011,      0.011,       0.011,       0.011,
  0.01126,    0.01126,     0.01126,     0.01126,
  0.01136,    0.01136,     0.01136,     0.01136,
  0.01143,    0.01143,     0.01143,     0.01143,
  0.01122,    0.01122,     0.01122,     0.01122,
  0.01128,    0.01128,     0.01128,     0.01128,
  0.01149,    0.01149,     0.01149,     0.01149,
  0.01136,    0.01136,     0.01136,     0.01136,
  0.01111,    0.01111,     0.01111,     0.01111,
  0.01058,    0.01058,     0.01058,     0.01058,
  0.01013,    0.01013,     0.01013,     0.01013,
  0.009901,   0.009901,    0.009901,    0.009901,
  0.009716,   0.009716,    0.009716,    0.009716,
  0.009694,   0.009694,    0.009694,    0.009694,
  0.009732,   0.009732,    0.009732,    0.009732,
  0.008705,   0.008705,    0.008705,    0.008705,
  0.007537,   0.007537,    0.007537,    0.007537,
  0.007408,   0.007408,    0.007408,    0.007408,
  0.007373,   0.007373,    0.007373,    0.007373,
  0.007362,   0.007362,    0.007362,    0.007362,
  0.007344,   0.007344,    0.007344,    0.007344,
  0.007407,   0.007407,    0.007407,    0.007407,
  0.007587,   0.007587,    0.007587,    0.007587,
  0.007691,   0.007691,    0.007691,    0.007691,
  0.007678,   0.007678,    0.007678,    0.007678,
  0.007778,   0.007778,    0.007778,    0.007778,
  0.008038,   0.008038,    0.008038,    0.008038,
  0.008366,   0.008366,    0.008366,    0.008366,
  0.008631,   0.008631,    0.008631,    0.008631,
  0.008756,   0.008756,    0.008756,    0.008756,
  0.00877,    0.00877,     0.00877,     0.00877,
  0.008614,   0.008614,    0.008614,    0.008614,
  0.008383,   0.008383,    0.008383,    0.008383,
  0.008058,   0.008058,    0.008058,    0.008058,
  0.007738,   0.007738,    0.007738,    0.007738,
  0.00755,    0.00755,     0.00755,     0.00755,
  0.007475,   0.007475,    0.007475,    0.007475,
  0.007295,   0.007295,    0.007295,    0.007295,
  0.006839,   0.006839,    0.006839,    0.006839,
  0.006433,   0.006433,    0.006433,    0.006433,
  0.006104,   0.006104,    0.006104,    0.006104,
  0.005726,   0.005726,    0.005726,    0.005726,
  0.005715,   0.005715,    0.005715,    0.005715,
  0.0075,     0.0075,      0.0075,      0.0075,
  0.00959,    0.00959,     0.00959,     0.00959,
  0.009977,   0.009977,    0.009977,    0.009977,
  0.009959,   0.009959,    0.009959,    0.009959,
  0.01005,    0.01005,     0.01005,     0.01005,
  0.009589,   0.009589,    0.009589,    0.009589,
  0.009311,   0.009311,    0.009311,    0.009311,
  0.009064,   0.009064,    0.009064,    0.009064,
  0.008888,   0.008888,    0.008888,    0.008888,
  0.009257,   0.009257,    0.009257,    0.009257,
  0.009141,   0.009141,    0.009141,    0.009141,
  0.008927,   0.008927,    0.008927,    0.008927,
  0.008992,   0.008992,    0.008992,    0.008992,
  0.009061,   0.009061,    0.009061,    0.009061,
  0.009031,   0.009031,    0.009031,    0.009031,
  0.009001,   0.009001,    0.009001,    0.009001,
  0.008995,   0.008995,    0.008995,    0.008995,
  0.009023,   0.009023,    0.009023,    0.009023,
  0.008945,   0.008945,    0.008945,    0.008945,
  0.008788,   0.008788,    0.008788,    0.008788,
  0.008709,   0.008709,    0.008709,    0.008709,
  0.008697,   0.008697,    0.008697,    0.008697,
  0.008753,   0.008753,    0.008753,    0.008753,
  0.008804,   0.008804,    0.008804,    0.008804,
  0.008854,   0.008854,    0.008854,    0.008854,
  0.00888,    0.00888,     0.00888,     0.00888,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.009111,   0.009111,    0.009111,    0.009111,
  0.009189,   0.009189,    0.009189,    0.009189,
  0.009242,   0.009242,    0.009242,    0.009242,
  0.009268,   0.009268,    0.009268,    0.009268,
  0.009263,   0.009263,    0.009263,    0.009263,
  0.009127,   0.009127,    0.009127,    0.009127,
  0.008812,   0.008812,    0.008812,    0.008812,
  0.008526,   0.008526,    0.008526,    0.008526,
  0.008403,   0.008403,    0.008403,    0.008403,
  0.008176,   0.008176,    0.008176,    0.008176,
  0.007808,   0.007808,    0.007808,    0.007808,
  0.007669,   0.007669,    0.007669,    0.007669,
  0.00825,    0.00825,     0.00825,     0.00825,
  0.008665,   0.008665,    0.008665,    0.008665,
  0.008148,   0.008148,    0.008148,    0.008148,
  0.007621,   0.007621,    0.007621,    0.007621,
  0.007399,   0.007399,    0.007399,    0.007399,
  0.007201,   0.007201,    0.007201,    0.007201,
  0.006942,   0.006942,    0.006942,    0.006942,
  0.006846,   0.006846,    0.006846,    0.006846,
  0.006626,   0.006626,    0.006626,    0.006626,
  0.006473,   0.006473,    0.006473,    0.006473,
  0.007178,   0.007178,    0.007178,    0.007178,
  0.008167,   0.008167,    0.008167,    0.008167,
  0.008591,   0.008591,    0.008591,    0.008591,
  0.008456,   0.008456,    0.008456,    0.008456,
  0.008322,   0.008322,    0.008322,    0.008322,
  0.008168,   0.008168,    0.008168,    0.008168,
  0.007867,   0.007867,    0.007867,    0.007867,
  0.007674,   0.007674,    0.007674,    0.007674,
  0.007681,   0.007681,    0.007681,    0.007681,
  0.00779,    0.00779,     0.00779,     0.00779,
  0.007912,   0.007912,    0.007912,    0.007912,
  0.008028,   0.008028,    0.008028,    0.008028,
  0.008052,   0.008052,    0.008052,    0.008052,
  0.008145,   0.008145,    0.008145,    0.008145,
  0.008328,   0.008328,    0.008328,    0.008328,
  0.008483,   0.008483,    0.008483,    0.008483,
  0.008597,   0.008597,    0.008597,    0.008597,
  0.008629,   0.008629,    0.008629,    0.008629,
  0.008629,   0.008629,    0.008629,    0.008629,
  0.008629,   0.008629,    0.008629,    0.008629,
  0.008629,   0.008629,    0.008629,    0.008629,
  0.008653,   0.008653,    0.008653,    0.008653,
  0.008678,   0.008678,    0.008678,    0.008678,
  0.008678,   0.008678,    0.008678,    0.008678,
  0.008678,   0.008678,    0.008678,    0.008678,
  0.008703,   0.008703,    0.008703,    0.008703,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008753,   0.008753,    0.008753,    0.008753,
  0.008804,   0.008804,    0.008804,    0.008804,
  0.00888,    0.00888,     0.00888,     0.00888,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.009111,   0.009111,    0.009111,    0.009111,
  0.009295,   0.009295,    0.009295,    0.009295,
  0.009428,   0.009428,    0.009428,    0.009428,
  0.009454,   0.009454,    0.009454,    0.009454,
  0.009508,   0.009508,    0.009508,    0.009508,
  0.009749,   0.009749,    0.009749,    0.009749,
  0.009915,   0.009915,    0.009915,    0.009915,
  0.009761,   0.009761,    0.009761,    0.009761,
  0.00956,    0.00956,     0.00956,     0.00956,
  0.009303,   0.009303,    0.009303,    0.009303,
  0.008992,   0.008992,    0.008992,    0.008992,
  0.008965,   0.008965,    0.008965,    0.008965,
  0.009062,   0.009062,    0.009062,    0.009062,
  0.009068,   0.009068,    0.009068,    0.009068,
  0.00907,    0.00907,     0.00907,     0.00907,
  0.008977,   0.008977,    0.008977,    0.008977,
  0.008977,   0.008977,    0.008977,    0.008977,
  0.009316,   0.009316,    0.009316,    0.009316,
  0.009622,   0.009622,    0.009622,    0.009622,
  0.00965,    0.00965,     0.00965,     0.00965,
  0.00968,    0.00968,     0.00968,     0.00968,
  0.009805,   0.009805,    0.009805,    0.009805,
  0.009838,   0.009838,    0.009838,    0.009838,
  0.009873,   0.009873,    0.009873,    0.009873,
  0.01001,    0.01001,     0.01001,     0.01001,
  0.01012,    0.01012,     0.01012,     0.01012,
  0.01012,    0.01012,     0.01012,     0.01012,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.009977,   0.009977,    0.009977,    0.009977,
  0.009921,   0.009921,    0.009921,    0.009921,
  0.009865,   0.009865,    0.009865,    0.009865,
  0.009837,   0.009837,    0.009837,    0.009837,
  0.009837,   0.009837,    0.009837,    0.009837,
  0.009865,   0.009865,    0.009865,    0.009865,
  0.009893,   0.009893,    0.009893,    0.009893,
  0.009921,   0.009921,    0.009921,    0.009921,
  0.009977,   0.009977,    0.009977,    0.009977,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.01015,    0.01015,     0.01015,     0.01015,
  0.0102,     0.0102,      0.0102,      0.0102,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.01026,    0.01026,     0.01026,     0.01026,
  0.01035,    0.01035,     0.01035,     0.01035,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01067,    0.01067,     0.01067,     0.01067,
  0.01079,    0.01079,     0.01079,     0.01079,
  0.01082,    0.01082,     0.01082,     0.01082,
  0.01085,    0.01085,     0.01085,     0.01085,
  0.01098,    0.01098,     0.01098,     0.01098,
  0.01088,    0.01088,     0.01088,     0.01088,
  0.0107,     0.0107,      0.0107,      0.0107,
  0.01053,    0.01053,     0.01053,     0.01053,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.009798,   0.009798,    0.009798,    0.009798,
  0.009453,   0.009453,    0.009453,    0.009453,
  0.009355,   0.009355,    0.009355,    0.009355,
  0.009158,   0.009158,    0.009158,    0.009158,
  0.008952,   0.008952,    0.008952,    0.008952,
  0.008894,   0.008894,    0.008894,    0.008894,
  0.00881,    0.00881,     0.00881,     0.00881,
  0.008616,   0.008616,    0.008616,    0.008616,
  0.008496,   0.008496,    0.008496,    0.008496,
  0.008451,   0.008451,    0.008451,    0.008451,
  0.008383,   0.008383,    0.008383,    0.008383,
  0.008366,   0.008366,    0.008366,    0.008366,
  0.008378,   0.008378,    0.008378,    0.008378,
  0.008315,   0.008315,    0.008315,    0.008315,
  0.008298,   0.008298,    0.008298,    0.008298,
  0.008482,   0.008482,    0.008482,    0.008482,
  0.00865,    0.00865,     0.00865,     0.00865,
  0.008646,   0.008646,    0.008646,    0.008646,
  0.008612,   0.008612,    0.008612,    0.008612,
  0.008735,   0.008735,    0.008735,    0.008735,
  0.008937,   0.008937,    0.008937,    0.008937,
  0.009138,   0.009138,    0.009138,    0.009138,
  0.009239,   0.009239,    0.009239,    0.009239,
  0.009124,   0.009124,    0.009124,    0.009124,
  0.009027,   0.009027,    0.009027,    0.009027,
  0.008976,   0.008976,    0.008976,    0.008976,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.009138,   0.009138,    0.009138,    0.009138,
  0.009189,   0.009189,    0.009189,    0.009189,
  0.009059,   0.009059,    0.009059,    0.009059,
  0.008855,   0.008855,    0.008855,    0.008855,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008804,   0.008804,    0.008804,    0.008804,
  0.00888,    0.00888,     0.00888,     0.00888,
  0.008854,   0.008854,    0.008854,    0.008854,
  0.008854,   0.008854,    0.008854,    0.008854,
  0.008905,   0.008905,    0.008905,    0.008905,
  0.009086,   0.009086,    0.009086,    0.009086,
  0.009375,   0.009375,    0.009375,    0.009375,
  0.009613,   0.009613,    0.009613,    0.009613,
  0.009667,   0.009667,    0.009667,    0.009667,
  0.009501,   0.009501,    0.009501,    0.009501,
  0.009285,   0.009285,    0.009285,    0.009285,
  0.009149,   0.009149,    0.009149,    0.009149,
  0.009114,   0.009114,    0.009114,    0.009114,
  0.008988,   0.008988,    0.008988,    0.008988,
  0.008867,   0.008867,    0.008867,    0.008867,
  0.00875,    0.00875,     0.00875,     0.00875,
  0.008601,   0.008601,    0.008601,    0.008601,
  0.008547,   0.008547,    0.008547,    0.008547,
  0.008419,   0.008419,    0.008419,    0.008419,
  0.008346,   0.008346,    0.008346,    0.008346,
  0.008364,   0.008364,    0.008364,    0.008364,
  0.008241,   0.008241,    0.008241,    0.008241,
  0.008276,   0.008276,    0.008276,    0.008276,
  0.00842,    0.00842,     0.00842,     0.00842,
  0.008445,   0.008445,    0.008445,    0.008445,
  0.008502,   0.008502,    0.008502,    0.008502,
  0.008625,   0.008625,    0.008625,    0.008625,
  0.008746,   0.008746,    0.008746,    0.008746,
  0.008828,   0.008828,    0.008828,    0.008828,
  0.008942,   0.008942,    0.008942,    0.008942,
  0.009091,   0.009091,    0.009091,    0.009091,
  0.009274,   0.009274,    0.009274,    0.009274,
  0.009366,   0.009366,    0.009366,    0.009366,
  0.009396,   0.009396,    0.009396,    0.009396,
  0.009396,   0.009396,    0.009396,    0.009396,
  0.009493,   0.009493,    0.009493,    0.009493,
  0.009687,   0.009687,    0.009687,    0.009687,
  0.009658,   0.009658,    0.009658,    0.009658,
  0.009503,   0.009503,    0.009503,    0.009503,
  0.009478,   0.009478,    0.009478,    0.009478,
  0.009521,   0.009521,    0.009521,    0.009521,
  0.009538,   0.009538,    0.009538,    0.009538,
  0.009523,   0.009523,    0.009523,    0.009523,
  0.009442,   0.009442,    0.009442,    0.009442,
  0.009235,   0.009235,    0.009235,    0.009235,
  0.008979,   0.008979,    0.008979,    0.008979,
  0.008789,   0.008789,    0.008789,    0.008789,
  0.008691,   0.008691,    0.008691,    0.008691,
  0.008643,   0.008643,    0.008643,    0.008643,
  0.008565,   0.008565,    0.008565,    0.008565,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.008623,   0.008623,    0.008623,    0.008623,
  0.008703,   0.008703,    0.008703,    0.008703,
  0.008791,   0.008791,    0.008791,    0.008791,
  0.008875,   0.008875,    0.008875,    0.008875,
  0.008884,   0.008884,    0.008884,    0.008884,
  0.008834,   0.008834,    0.008834,    0.008834,
  0.008781,   0.008781,    0.008781,    0.008781,
  0.008738,   0.008738,    0.008738,    0.008738,
  0.008548,   0.008548,    0.008548,    0.008548,
  0.008181,   0.008181,    0.008181,    0.008181,
  0.007843,   0.007843,    0.007843,    0.007843,
  0.0077,     0.0077,      0.0077,      0.0077,
  0.007759,   0.007759,    0.007759,    0.007759,
  0.007693,   0.007693,    0.007693,    0.007693,
  0.007669,   0.007669,    0.007669,    0.007669,
  0.007782,   0.007782,    0.007782,    0.007782,
  0.007798,   0.007798,    0.007798,    0.007798,
  0.007892,   0.007892,    0.007892,    0.007892,
  0.007982,   0.007982,    0.007982,    0.007982,
  0.008028,   0.008028,    0.008028,    0.008028,
  0.007965,   0.007965,    0.007965,    0.007965,
  0.007913,   0.007913,    0.007913,    0.007913,
  0.007971,   0.007971,    0.007971,    0.007971,
  0.008002,   0.008002,    0.008002,    0.008002,
  0.008034,   0.008034,    0.008034,    0.008034,
  0.007998,   0.007998,    0.007998,    0.007998,
  0.007988,   0.007988,    0.007988,    0.007988,
  0.007857,   0.007857,    0.007857,    0.007857,
  0.007759,   0.007759,    0.007759,    0.007759,
  0.007924,   0.007924,    0.007924,    0.007924,
  0.008108,   0.008108,    0.008108,    0.008108,
  0.008252,   0.008252,    0.008252,    0.008252,
  0.00832,    0.00832,     0.00832,     0.00832,
  0.008267,   0.008267,    0.008267,    0.008267,
  0.00824,    0.00824,     0.00824,     0.00824,
  0.008236,   0.008236,    0.008236,    0.008236,
  0.008161,   0.008161,    0.008161,    0.008161,
  0.008061,   0.008061,    0.008061,    0.008061,
  0.008,      0.008,       0.008,       0.008,
  0.007973,   0.007973,    0.007973,    0.007973,
  0.007954,   0.007954,    0.007954,    0.007954,
  0.007922,   0.007922,    0.007922,    0.007922,
  0.007847,   0.007847,    0.007847,    0.007847,
  0.007785,   0.007785,    0.007785,    0.007785,
  0.007747,   0.007747,    0.007747,    0.007747,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007394,   0.007394,    0.007394,    0.007394,
  0.007218,   0.007218,    0.007218,    0.007218,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007304,   0.007304,    0.007304,    0.007304,
  0.007446,   0.007446,    0.007446,    0.007446,
  0.007769,   0.007769,    0.007769,    0.007769,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008117,   0.008117,    0.008117,    0.008117,
  0.007975,   0.007975,    0.007975,    0.007975,
  0.007866,   0.007866,    0.007866,    0.007866,
  0.007848,   0.007848,    0.007848,    0.007848,
  0.007799,   0.007799,    0.007799,    0.007799,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007609,   0.007609,    0.007609,    0.007609,
  0.007441,   0.007441,    0.007441,    0.007441,
  0.007256,   0.007256,    0.007256,    0.007256,
  0.007116,   0.007116,    0.007116,    0.007116,
  0.006942,   0.006942,    0.006942,    0.006942,
  0.006841,   0.006841,    0.006841,    0.006841,
  0.006787,   0.006787,    0.006787,    0.006787,
  0.006879,   0.006879,    0.006879,    0.006879,
  0.00704,    0.00704,     0.00704,     0.00704,
  0.006734,   0.006734,    0.006734,    0.006734,
  0.006662,   0.006662,    0.006662,    0.006662,
  0.006751,   0.006751,    0.006751,    0.006751,
  0.006292,   0.006292,    0.006292,    0.006292,
  0.006166,   0.006166,    0.006166,    0.006166,
  0.006345,   0.006345,    0.006345,    0.006345,
  0.006931,   0.006931,    0.006931,    0.006931,
  0.007406,   0.007406,    0.007406,    0.007406,
  0.0076,     0.0076,      0.0076,      0.0076,
  0.008065,   0.008065,    0.008065,    0.008065,
  0.00841,    0.00841,     0.00841,     0.00841,
  0.008519,   0.008519,    0.008519,    0.008519,
  0.00847,    0.00847,     0.00847,     0.00847,
  0.00846,    0.00846,     0.00846,     0.00846,
  0.008611,   0.008611,    0.008611,    0.008611,
  0.008924,   0.008924,    0.008924,    0.008924,
  0.009302,   0.009302,    0.009302,    0.009302,
  0.009525,   0.009525,    0.009525,    0.009525,
  0.009528,   0.009528,    0.009528,    0.009528,
  0.009438,   0.009438,    0.009438,    0.009438,
  0.009316,   0.009316,    0.009316,    0.009316,
  0.00916,    0.00916,     0.00916,     0.00916,
  0.009004,   0.009004,    0.009004,    0.009004,
  0.008883,   0.008883,    0.008883,    0.008883,
  0.008796,   0.008796,    0.008796,    0.008796,
  0.008711,   0.008711,    0.008711,    0.008711,
  0.008633,   0.008633,    0.008633,    0.008633,
  0.008619,   0.008619,    0.008619,    0.008619,
  0.008601,   0.008601,    0.008601,    0.008601,
  0.008595,   0.008595,    0.008595,    0.008595,
  0.008626,   0.008626,    0.008626,    0.008626,
  0.008626,   0.008626,    0.008626,    0.008626,
  0.00858,    0.00858,     0.00858,     0.00858,
  0.008558,   0.008558,    0.008558,    0.008558,
  0.008594,   0.008594,    0.008594,    0.008594,
  0.008567,   0.008567,    0.008567,    0.008567,
  0.008528,   0.008528,    0.008528,    0.008528,
  0.008367,   0.008367,    0.008367,    0.008367,
  0.008207,   0.008207,    0.008207,    0.008207,
  0.007891,   0.007891,    0.007891,    0.007891,
  0.007353,   0.007353,    0.007353,    0.007353,
  0.007053,   0.007053,    0.007053,    0.007053,
  0.006852,   0.006852,    0.006852,    0.006852,
  0.006624,   0.006624,    0.006624,    0.006624,
  0.006537,   0.006537,    0.006537,    0.006537,
  0.0065,     0.0065,      0.0065,      0.0065,
  0.006397,   0.006397,    0.006397,    0.006397,
  0.006187,   0.006187,    0.006187,    0.006187,
  0.006078,   0.006078,    0.006078,    0.006078,
  0.006176,   0.006176,    0.006176,    0.006176,
  0.006064,   0.006064,    0.006064,    0.006064,
  0.005907,   0.005907,    0.005907,    0.005907,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.006096,   0.006096,    0.006096,    0.006096,
  0.006303,   0.006303,    0.006303,    0.006303,
  0.006604,   0.006604,    0.006604,    0.006604,
  0.006914,   0.006914,    0.006914,    0.006914,
  0.007256,   0.007256,    0.007256,    0.007256,
  0.007602,   0.007602,    0.007602,    0.007602,
  0.00782,    0.00782,     0.00782,     0.00782,
  0.00793,    0.00793,     0.00793,     0.00793,
  0.008028,   0.008028,    0.008028,    0.008028,
  0.008114,   0.008114,    0.008114,    0.008114,
  0.008165,   0.008165,    0.008165,    0.008165,
  0.008203,   0.008203,    0.008203,    0.008203,
  0.008303,   0.008303,    0.008303,    0.008303,
  0.008441,   0.008441,    0.008441,    0.008441,
  0.008491,   0.008491,    0.008491,    0.008491,
  0.008546,   0.008546,    0.008546,    0.008546,
  0.008609,   0.008609,    0.008609,    0.008609,
  0.008642,   0.008642,    0.008642,    0.008642,
  0.008709,   0.008709,    0.008709,    0.008709,
  0.00878,    0.00878,     0.00878,     0.00878,
  0.008856,   0.008856,    0.008856,    0.008856,
  0.008966,   0.008966,    0.008966,    0.008966,
  0.009102,   0.009102,    0.009102,    0.009102,
  0.009228,   0.009228,    0.009228,    0.009228,
  0.009338,   0.009338,    0.009338,    0.009338,
  0.009471,   0.009471,    0.009471,    0.009471,
  0.009491,   0.009491,    0.009491,    0.009491,
  0.009432,   0.009432,    0.009432,    0.009432,
  0.009453,   0.009453,    0.009453,    0.009453,
  0.009478,   0.009478,    0.009478,    0.009478,
  0.009413,   0.009413,    0.009413,    0.009413,
  0.00928,    0.00928,     0.00928,     0.00928,
  0.009123,   0.009123,    0.009123,    0.009123,
  0.008834,   0.008834,    0.008834,    0.008834,
  0.008365,   0.008365,    0.008365,    0.008365,
  0.007721,   0.007721,    0.007721,    0.007721,
  0.007257,   0.007257,    0.007257,    0.007257,
  0.007103,   0.007103,    0.007103,    0.007103,
  0.007185,   0.007185,    0.007185,    0.007185,
  0.007135,   0.007135,    0.007135,    0.007135,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.007181,   0.007181,    0.007181,    0.007181,
  0.007063,   0.007063,    0.007063,    0.007063,
  0.007029,   0.007029,    0.007029,    0.007029,
  0.007059,   0.007059,    0.007059,    0.007059,
  0.007122,   0.007122,    0.007122,    0.007122,
  0.00725,    0.00725,     0.00725,     0.00725,
  0.007364,   0.007364,    0.007364,    0.007364,
  0.00737,    0.00737,     0.00737,     0.00737,
  0.00736,    0.00736,     0.00736,     0.00736,
  0.007483,   0.007483,    0.007483,    0.007483,
  0.007599,   0.007599,    0.007599,    0.007599,
  0.007636,   0.007636,    0.007636,    0.007636,
  0.007558,   0.007558,    0.007558,    0.007558,
  0.007281,   0.007281,    0.007281,    0.007281,
  0.006918,   0.006918,    0.006918,    0.006918,
  0.006752,   0.006752,    0.006752,    0.006752,
  0.006759,   0.006759,    0.006759,    0.006759,
  0.006827,   0.006827,    0.006827,    0.006827,
  0.006901,   0.006901,    0.006901,    0.006901,
  0.006969,   0.006969,    0.006969,    0.006969,
  0.007158,   0.007158,    0.007158,    0.007158,
  0.007391,   0.007391,    0.007391,    0.007391,
  0.007573,   0.007573,    0.007573,    0.007573,
  0.007728,   0.007728,    0.007728,    0.007728,
  0.007822,   0.007822,    0.007822,    0.007822,
  0.007884,   0.007884,    0.007884,    0.007884,
  0.007947,   0.007947,    0.007947,    0.007947,
  0.008011,   0.008011,    0.008011,    0.008011,
  0.008107,   0.008107,    0.008107,    0.008107,
  0.008209,   0.008209,    0.008209,    0.008209,
  0.008312,   0.008312,    0.008312,    0.008312,
  0.008472,   0.008472,    0.008472,    0.008472,
  0.008619,   0.008619,    0.008619,    0.008619,
  0.008642,   0.008642,    0.008642,    0.008642,
  0.008684,   0.008684,    0.008684,    0.008684,
  0.008763,   0.008763,    0.008763,    0.008763,
  0.008739,   0.008739,    0.008739,    0.008739,
  0.008627,   0.008627,    0.008627,    0.008627,
  0.00841,    0.00841,     0.00841,     0.00841,
  0.008179,   0.008179,    0.008179,    0.008179,
  0.007689,   0.007689,    0.007689,    0.007689,
  0.007176,   0.007176,    0.007176,    0.007176,
  0.006926,   0.006926,    0.006926,    0.006926,
  0.006511,   0.006511,    0.006511,    0.006511,
  0.006097,   0.006097,    0.006097,    0.006097,
  0.005765,   0.005765,    0.005765,    0.005765,
  0.005639,   0.005639,    0.005639,    0.005639,
  0.005702,   0.005702,    0.005702,    0.005702,
  0.005674,   0.005674,    0.005674,    0.005674,
  0.005615,   0.005615,    0.005615,    0.005615,
  0.005487,   0.005487,    0.005487,    0.005487,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.00516,    0.00516,     0.00516,     0.00516,
  0.005472,   0.005472,    0.005472,    0.005472,
  0.005717,   0.005717,    0.005717,    0.005717,
  0.005812,   0.005812,    0.005812,    0.005812,
  0.006127,   0.006127,    0.006127,    0.006127,
  0.006638,   0.006638,    0.006638,    0.006638,
  0.007264,   0.007264,    0.007264,    0.007264,
  0.007739,   0.007739,    0.007739,    0.007739,
  0.00817,    0.00817,     0.00817,     0.00817,
  0.008543,   0.008543,    0.008543,    0.008543,
  0.008667,   0.008667,    0.008667,    0.008667,
  0.008766,   0.008766,    0.008766,    0.008766,
  0.008885,   0.008885,    0.008885,    0.008885,
  0.008854,   0.008854,    0.008854,    0.008854,
  0.008868,   0.008868,    0.008868,    0.008868,
  0.008883,   0.008883,    0.008883,    0.008883,
  0.008817,   0.008817,    0.008817,    0.008817,
  0.008843,   0.008843,    0.008843,    0.008843,
  0.00893,    0.00893,     0.00893,     0.00893,
  0.008944,   0.008944,    0.008944,    0.008944,
  0.008994,   0.008994,    0.008994,    0.008994,
  0.00899,    0.00899,     0.00899,     0.00899,
  0.008924,   0.008924,    0.008924,    0.008924,
  0.008988,   0.008988,    0.008988,    0.008988,
  0.009119,   0.009119,    0.009119,    0.009119,
  0.009192,   0.009192,    0.009192,    0.009192,
  0.009196,   0.009196,    0.009196,    0.009196,
  0.009253,   0.009253,    0.009253,    0.009253,
  0.009338,   0.009338,    0.009338,    0.009338,
  0.00942,    0.00942,     0.00942,     0.00942,
  0.009379,   0.009379,    0.009379,    0.009379,
  0.009218,   0.009218,    0.009218,    0.009218,
  0.008998,   0.008998,    0.008998,    0.008998,
  0.008544,   0.008544,    0.008544,    0.008544,
  0.007961,   0.007961,    0.007961,    0.007961,
  0.007233,   0.007233,    0.007233,    0.007233,
  0.006347,   0.006347,    0.006347,    0.006347,
  0.005927,   0.005927,    0.005927,    0.005927,
  0.005834,   0.005834,    0.005834,    0.005834,
  0.005624,   0.005624,    0.005624,    0.005624,
  0.005876,   0.005876,    0.005876,    0.005876,
  0.006083,   0.006083,    0.006083,    0.006083,
  0.005959,   0.005959,    0.005959,    0.005959,
  0.00561,    0.00561,     0.00561,     0.00561,
  0.005188,   0.005188,    0.005188,    0.005188,
  0.005188,   0.005188,    0.005188,    0.005188,
  0.005268,   0.005268,    0.005268,    0.005268,
  0.005305,   0.005305,    0.005305,    0.005305,
  0.005388,   0.005388,    0.005388,    0.005388,
  0.006431,   0.006431,    0.006431,    0.006431,
  0.007194,   0.007194,    0.007194,    0.007194,
  0.007045,   0.007045,    0.007045,    0.007045,
  0.0072,     0.0072,      0.0072,      0.0072,
  0.007423,   0.007423,    0.007423,    0.007423,
  0.007935,   0.007935,    0.007935,    0.007935,
  0.008676,   0.008676,    0.008676,    0.008676,
  0.008662,   0.008662,    0.008662,    0.008662,
  0.008476,   0.008476,    0.008476,    0.008476,
  0.008597,   0.008597,    0.008597,    0.008597,
  0.008496,   0.008496,    0.008496,    0.008496,
  0.008662,   0.008662,    0.008662,    0.008662,
  0.009029,   0.009029,    0.009029,    0.009029,
  0.009243,   0.009243,    0.009243,    0.009243,
  0.009284,   0.009284,    0.009284,    0.009284,
  0.009182,   0.009182,    0.009182,    0.009182,
  0.009078,   0.009078,    0.009078,    0.009078,
  0.009067,   0.009067,    0.009067,    0.009067,
  0.009002,   0.009002,    0.009002,    0.009002,
  0.008937,   0.008937,    0.008937,    0.008937,
  0.008701,   0.008701,    0.008701,    0.008701,
  0.008421,   0.008421,    0.008421,    0.008421,
  0.008372,   0.008372,    0.008372,    0.008372,
  0.008335,   0.008335,    0.008335,    0.008335,
  0.008266,   0.008266,    0.008266,    0.008266,
  0.008175,   0.008175,    0.008175,    0.008175,
  0.008239,   0.008239,    0.008239,    0.008239,
  0.008642,   0.008642,    0.008642,    0.008642,
  0.009188,   0.009188,    0.009188,    0.009188,
  0.009509,   0.009509,    0.009509,    0.009509,
  0.009337,   0.009337,    0.009337,    0.009337,
  0.008925,   0.008925,    0.008925,    0.008925,
  0.008588,   0.008588,    0.008588,    0.008588,
  0.008165,   0.008165,    0.008165,    0.008165,
  0.007223,   0.007223,    0.007223,    0.007223,
  0.006022,   0.006022,    0.006022,    0.006022,
  0.005228,   0.005228,    0.005228,    0.005228,
  0.004572,   0.004572,    0.004572,    0.004572,
  0.004259,   0.004259,    0.004259,    0.004259,
  0.004355,   0.004355,    0.004355,    0.004355,
  0.004324,   0.004324,    0.004324,    0.004324,
  0.004333,   0.004333,    0.004333,    0.004333,
  0.004305,   0.004305,    0.004305,    0.004305,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004422,   0.004422,    0.004422,    0.004422,
  0.004598,   0.004598,    0.004598,    0.004598,
  0.004264,   0.004264,    0.004264,    0.004264,
  0.004066,   0.004066,    0.004066,    0.004066,
  0.004044,   0.004044,    0.004044,    0.004044,
  0.004,      0.004,       0.004,       0.004,
  0.004385,   0.004385,    0.004385,    0.004385,
  0.004982,   0.004982,    0.004982,    0.004982,
  0.005549,   0.005549,    0.005549,    0.005549,
  0.006054,   0.006054,    0.006054,    0.006054,
  0.006447,   0.006447,    0.006447,    0.006447,
  0.006751,   0.006751,    0.006751,    0.006751,
  0.006979,   0.006979,    0.006979,    0.006979,
  0.007082,   0.007082,    0.007082,    0.007082,
  0.007101,   0.007101,    0.007101,    0.007101,
  0.007028,   0.007028,    0.007028,    0.007028,
  0.007065,   0.007065,    0.007065,    0.007065,
  0.007242,   0.007242,    0.007242,    0.007242,
  0.007208,   0.007208,    0.007208,    0.007208,
  0.007098,   0.007098,    0.007098,    0.007098,
  0.007202,   0.007202,    0.007202,    0.007202,
  0.007316,   0.007316,    0.007316,    0.007316,
  0.007356,   0.007356,    0.007356,    0.007356,
  0.0074,     0.0074,      0.0074,      0.0074,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007683,   0.007683,    0.007683,    0.007683,
  0.007811,   0.007811,    0.007811,    0.007811,
  0.007863,   0.007863,    0.007863,    0.007863,
  0.00786,    0.00786,     0.00786,     0.00786,
  0.007859,   0.007859,    0.007859,    0.007859,
  0.007831,   0.007831,    0.007831,    0.007831,
  0.007752,   0.007752,    0.007752,    0.007752,
  0.007663,   0.007663,    0.007663,    0.007663,
  0.007414,   0.007414,    0.007414,    0.007414,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.006912,   0.006912,    0.006912,    0.006912,
  0.006857,   0.006857,    0.006857,    0.006857,
  0.006823,   0.006823,    0.006823,    0.006823,
  0.006671,   0.006671,    0.006671,    0.006671,
  0.006357,   0.006357,    0.006357,    0.006357,
  0.005752,   0.005752,    0.005752,    0.005752,
  0.005134,   0.005134,    0.005134,    0.005134,
  0.004714,   0.004714,    0.004714,    0.004714,
  0.004524,   0.004524,    0.004524,    0.004524,
  0.004453,   0.004453,    0.004453,    0.004453,
  0.004205,   0.004205,    0.004205,    0.004205,
  0.004048,   0.004048,    0.004048,    0.004048,
  0.003833,   0.003833,    0.003833,    0.003833,
  0.003559,   0.003559,    0.003559,    0.003559,
  0.003171,   0.003171,    0.003171,    0.003171,
  0.002777,   0.002777,    0.002777,    0.002777,
  0.002541,   0.002541,    0.002541,    0.002541,
  0.002337,   0.002337,    0.002337,    0.002337,
  0.002455,   0.002455,    0.002455,    0.002455,
  0.002912,   0.002912,    0.002912,    0.002912,
  0.00356,    0.00356,     0.00356,     0.00356,
  0.004127,   0.004127,    0.004127,    0.004127,
  0.004692,   0.004692,    0.004692,    0.004692,
  0.005267,   0.005267,    0.005267,    0.005267,
  0.00573,    0.00573,     0.00573,     0.00573,
  0.00603,    0.00603,     0.00603,     0.00603,
  0.006261,   0.006261,    0.006261,    0.006261,
  0.00645,    0.00645,     0.00645,     0.00645,
  0.006548,   0.006548,    0.006548,    0.006548,
  0.006703,   0.006703,    0.006703,    0.006703,
  0.006878,   0.006878,    0.006878,    0.006878,
  0.006934,   0.006934,    0.006934,    0.006934,
  0.006867,   0.006867,    0.006867,    0.006867,
  0.006772,   0.006772,    0.006772,    0.006772,
  0.006797,   0.006797,    0.006797,    0.006797,
  0.00689,    0.00689,     0.00689,     0.00689,
  0.007001,   0.007001,    0.007001,    0.007001,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007153,   0.007153,    0.007153,    0.007153,
  0.007198,   0.007198,    0.007198,    0.007198,
  0.007185,   0.007185,    0.007185,    0.007185,
  0.007255,   0.007255,    0.007255,    0.007255,
  0.007484,   0.007484,    0.007484,    0.007484,
  0.007698,   0.007698,    0.007698,    0.007698,
  0.007873,   0.007873,    0.007873,    0.007873,
  0.007825,   0.007825,    0.007825,    0.007825,
  0.007448,   0.007448,    0.007448,    0.007448,
  0.00695,    0.00695,     0.00695,     0.00695,
  0.006445,   0.006445,    0.006445,    0.006445,
  0.006055,   0.006055,    0.006055,    0.006055,
  0.005819,   0.005819,    0.005819,    0.005819,
  0.005661,   0.005661,    0.005661,    0.005661,
  0.005613,   0.005613,    0.005613,    0.005613,
  0.005578,   0.005578,    0.005578,    0.005578,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.004257,   0.004257,    0.004257,    0.004257,
  0.003569,   0.003569,    0.003569,    0.003569,
  0.003216,   0.003216,    0.003216,    0.003216,
  0.003144,   0.003144,    0.003144,    0.003144,
  0.003306,   0.003306,    0.003306,    0.003306,
  0.003195,   0.003195,    0.003195,    0.003195,
  0.002919,   0.002919,    0.002919,    0.002919,
  0.002974,   0.002974,    0.002974,    0.002974,
  0.003029,   0.003029,    0.003029,    0.003029,
  0.003135,   0.003135,    0.003135,    0.003135,
  0.003578,   0.003578,    0.003578,    0.003578,
  0.00384,    0.00384,     0.00384,     0.00384,
  0.003725,   0.003725,    0.003725,    0.003725,
  0.003744,   0.003744,    0.003744,    0.003744,
  0.004187,   0.004187,    0.004187,    0.004187,
  0.004849,   0.004849,    0.004849,    0.004849,
  0.005729,   0.005729,    0.005729,    0.005729,
  0.006535,   0.006535,    0.006535,    0.006535,
  0.006774,   0.006774,    0.006774,    0.006774,
  0.006882,   0.006882,    0.006882,    0.006882,
  0.007115,   0.007115,    0.007115,    0.007115,
  0.007232,   0.007232,    0.007232,    0.007232,
  0.007298,   0.007298,    0.007298,    0.007298,
  0.007376,   0.007376,    0.007376,    0.007376,
  0.007325,   0.007325,    0.007325,    0.007325,
  0.007327,   0.007327,    0.007327,    0.007327,
  0.007463,   0.007463,    0.007463,    0.007463,
  0.007469,   0.007469,    0.007469,    0.007469,
  0.00739,    0.00739,     0.00739,     0.00739,
  0.007296,   0.007296,    0.007296,    0.007296,
  0.007359,   0.007359,    0.007359,    0.007359,
  0.007581,   0.007581,    0.007581,    0.007581,
  0.007727,   0.007727,    0.007727,    0.007727,
  0.007821,   0.007821,    0.007821,    0.007821,
  0.007853,   0.007853,    0.007853,    0.007853,
  0.007853,   0.007853,    0.007853,    0.007853,
  0.007915,   0.007915,    0.007915,    0.007915,
  0.00801,    0.00801,     0.00801,     0.00801,
  0.008107,   0.008107,    0.008107,    0.008107,
  0.008139,   0.008139,    0.008139,    0.008139,
  0.00792,    0.00792,     0.00792,     0.00792,
  0.007561,   0.007561,    0.007561,    0.007561,
  0.007232,   0.007232,    0.007232,    0.007232,
  0.007108,   0.007108,    0.007108,    0.007108,
  0.007079,   0.007079,    0.007079,    0.007079,
  0.006718,   0.006718,    0.006718,    0.006718,
  0.005388,   0.005388,    0.005388,    0.005388,
  0.003678,   0.003678,    0.003678,    0.003678,
  0.002559,   0.002559,    0.002559,    0.002559,
  0.002033,   0.002033,    0.002033,    0.002033,
  0.002076,   0.002076,    0.002076,    0.002076,
  0.00224,    0.00224,     0.00224,     0.00224,
  0.002234,   0.002234,    0.002234,    0.002234,
  0.002486,   0.002486,    0.002486,    0.002486,
  0.002807,   0.002807,    0.002807,    0.002807,
  0.00333,    0.00333,     0.00333,     0.00333,
  0.004035,   0.004035,    0.004035,    0.004035,
  0.004585,   0.004585,    0.004585,    0.004585,
  0.005156,   0.005156,    0.005156,    0.005156,
  0.005622,   0.005622,    0.005622,    0.005622,
  0.0061,     0.0061,      0.0061,      0.0061,
  0.006697,   0.006697,    0.006697,    0.006697,
  0.007085,   0.007085,    0.007085,    0.007085,
  0.00735,    0.00735,     0.00735,     0.00735,
  0.008099,   0.008099,    0.008099,    0.008099,
  0.008907,   0.008907,    0.008907,    0.008907,
  0.009212,   0.009212,    0.009212,    0.009212,
  0.009269,   0.009269,    0.009269,    0.009269,
  0.009521,   0.009521,    0.009521,    0.009521,
  0.009941,   0.009941,    0.009941,    0.009941,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01054,    0.01054,     0.01054,     0.01054,
  0.01064,    0.01064,     0.01064,     0.01064,
  0.01072,    0.01072,     0.01072,     0.01072,
  0.01069,    0.01069,     0.01069,     0.01069,
  0.0106,     0.0106,      0.0106,      0.0106,
  0.01057,    0.01057,     0.01057,     0.01057,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01034,    0.01034,     0.01034,     0.01034,
  0.01017,    0.01017,     0.01017,     0.01017,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.009921,   0.009921,    0.009921,    0.009921,
  0.009782,   0.009782,    0.009782,    0.009782,
  0.009782,   0.009782,    0.009782,    0.009782,
  0.01001,    0.01001,     0.01001,     0.01001,
  0.0102,     0.0102,      0.0102,      0.0102,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01053,    0.01053,     0.01053,     0.01053,
  0.01067,    0.01067,     0.01067,     0.01067,
  0.01082,    0.01082,     0.01082,     0.01082,
  0.0111,     0.0111,      0.0111,      0.0111,
  0.01132,    0.01132,     0.01132,     0.01132,
  0.01123,    0.01123,     0.01123,     0.01123,
  0.01095,    0.01095,     0.01095,     0.01095,
  0.01087,    0.01087,     0.01087,     0.01087,
  0.01089,    0.01089,     0.01089,     0.01089,
  0.01083,    0.01083,     0.01083,     0.01083,
  0.01077,    0.01077,     0.01077,     0.01077,
  0.0107,     0.0107,      0.0107,      0.0107,
  0.01063,    0.01063,     0.01063,     0.01063,
  0.01062,    0.01062,     0.01062,     0.01062,
  0.01063,    0.01063,     0.01063,     0.01063,
  0.01054,    0.01054,     0.01054,     0.01054,
  0.01047,    0.01047,     0.01047,     0.01047,
  0.01028,    0.01028,     0.01028,     0.01028,
  0.00992,    0.00992,     0.00992,     0.00992,
  0.009735,   0.009735,    0.009735,    0.009735,
  0.009599,   0.009599,    0.009599,    0.009599,
  0.009596,   0.009596,    0.009596,    0.009596,
  0.009787,   0.009787,    0.009787,    0.009787,
  0.01002,    0.01002,     0.01002,     0.01002,
  0.01024,    0.01024,     0.01024,     0.01024,
  0.01036,    0.01036,     0.01036,     0.01036,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01022,    0.01022,     0.01022,     0.01022,
  0.01022,    0.01022,     0.01022,     0.01022,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.01022,    0.01022,     0.01022,     0.01022,
  0.01022,    0.01022,     0.01022,     0.01022,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.01018,    0.01018,     0.01018,     0.01018,
  0.01005,    0.01005,     0.01005,     0.01005,
  0.009862,   0.009862,    0.009862,    0.009862,
  0.009754,   0.009754,    0.009754,    0.009754,
  0.009644,   0.009644,    0.009644,    0.009644,
  0.009508,   0.009508,    0.009508,    0.009508,
  0.009401,   0.009401,    0.009401,    0.009401,
  0.009374,   0.009374,    0.009374,    0.009374,
  0.009428,   0.009428,    0.009428,    0.009428,
  0.009508,   0.009508,    0.009508,    0.009508,
  0.009617,   0.009617,    0.009617,    0.009617,
  0.009838,   0.009838,    0.009838,    0.009838,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01067,    0.01067,     0.01067,     0.01067,
  0.01056,    0.01056,     0.01056,     0.01056,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.009871,   0.009871,    0.009871,    0.009871,
  0.009631,   0.009631,    0.009631,    0.009631,
  0.009363,   0.009363,    0.009363,    0.009363,
  0.009134,   0.009134,    0.009134,    0.009134,
  0.008947,   0.008947,    0.008947,    0.008947,
  0.008657,   0.008657,    0.008657,    0.008657,
  0.008047,   0.008047,    0.008047,    0.008047,
  0.00776,    0.00776,     0.00776,     0.00776,
  0.007877,   0.007877,    0.007877,    0.007877,
  0.007792,   0.007792,    0.007792,    0.007792,
  0.007556,   0.007556,    0.007556,    0.007556,
  0.007333,   0.007333,    0.007333,    0.007333,
  0.007552,   0.007552,    0.007552,    0.007552,
  0.008311,   0.008311,    0.008311,    0.008311,
  0.008805,   0.008805,    0.008805,    0.008805,
  0.008744,   0.008744,    0.008744,    0.008744,
  0.008627,   0.008627,    0.008627,    0.008627,
  0.008612,   0.008612,    0.008612,    0.008612,
  0.008718,   0.008718,    0.008718,    0.008718,
  0.009019,   0.009019,    0.009019,    0.009019,
  0.009342,   0.009342,    0.009342,    0.009342,
  0.009376,   0.009376,    0.009376,    0.009376,
  0.009428,   0.009428,    0.009428,    0.009428,
  0.009682,   0.009682,    0.009682,    0.009682,
  0.009818,   0.009818,    0.009818,    0.009818,
  0.009706,   0.009706,    0.009706,    0.009706,
  0.009753,   0.009753,    0.009753,    0.009753,
  0.009892,   0.009892,    0.009892,    0.009892,
  0.00982,    0.00982,     0.00982,     0.00982,
  0.009833,   0.009833,    0.009833,    0.009833,
  0.009782,   0.009782,    0.009782,    0.009782,
  0.00943,    0.00943,     0.00943,     0.00943,
  0.008959,   0.008959,    0.008959,    0.008959,
  0.008532,   0.008532,    0.008532,    0.008532,
  0.008633,   0.008633,    0.008633,    0.008633,
  0.008804,   0.008804,    0.008804,    0.008804,
  0.008388,   0.008388,    0.008388,    0.008388,
  0.008241,   0.008241,    0.008241,    0.008241,
  0.008432,   0.008432,    0.008432,    0.008432,
  0.008384,   0.008384,    0.008384,    0.008384,
  0.008533,   0.008533,    0.008533,    0.008533,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008754,   0.008754,    0.008754,    0.008754,
  0.009361,   0.009361,    0.009361,    0.009361,
  0.01036,    0.01036,     0.01036,     0.01036,
  0.01098,    0.01098,     0.01098,     0.01098,
  0.01098,    0.01098,     0.01098,     0.01098,
  0.01033,    0.01033,     0.01033,     0.01033,
  0.009583,   0.009583,    0.009583,    0.009583,
  0.009023,   0.009023,    0.009023,    0.009023,
  0.008736,   0.008736,    0.008736,    0.008736,
  0.00844,    0.00844,     0.00844,     0.00844,
  0.007913,   0.007913,    0.007913,    0.007913,
  0.007617,   0.007617,    0.007617,    0.007617,
  0.007351,   0.007351,    0.007351,    0.007351,
  0.007269,   0.007269,    0.007269,    0.007269,
  0.00713,    0.00713,     0.00713,     0.00713,
  0.007019,   0.007019,    0.007019,    0.007019,
  0.007291,   0.007291,    0.007291,    0.007291,
  0.007512,   0.007512,    0.007512,    0.007512,
  0.007627,   0.007627,    0.007627,    0.007627,
  0.007469,   0.007469,    0.007469,    0.007469,
  0.007291,   0.007291,    0.007291,    0.007291,
  0.007722,   0.007722,    0.007722,    0.007722,
  0.008432,   0.008432,    0.008432,    0.008432,
  0.008856,   0.008856,    0.008856,    0.008856,
  0.009043,   0.009043,    0.009043,    0.009043,
  0.009255,   0.009255,    0.009255,    0.009255,
  0.009548,   0.009548,    0.009548,    0.009548,
  0.009779,   0.009779,    0.009779,    0.009779,
  0.009915,   0.009915,    0.009915,    0.009915,
  0.01002,    0.01002,     0.01002,     0.01002,
  0.0101,     0.0101,      0.0101,      0.0101,
  0.01013,    0.01013,     0.01013,     0.01013,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.009964,   0.009964,    0.009964,    0.009964,
  0.009934,   0.009934,    0.009934,    0.009934,
  0.00991,    0.00991,     0.00991,     0.00991,
  0.009891,   0.009891,    0.009891,    0.009891,
  0.009867,   0.009867,    0.009867,    0.009867,
  0.009811,   0.009811,    0.009811,    0.009811,
  0.009735,   0.009735,    0.009735,    0.009735,
  0.009655,   0.009655,    0.009655,    0.009655,
  0.009582,   0.009582,    0.009582,    0.009582,
  0.009514,   0.009514,    0.009514,    0.009514,
  0.009414,   0.009414,    0.009414,    0.009414,
  0.009311,   0.009311,    0.009311,    0.009311,
  0.00929,    0.00929,     0.00929,     0.00929,
  0.009424,   0.009424,    0.009424,    0.009424,
  0.00971,    0.00971,     0.00971,     0.00971,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.01019,    0.01019,     0.01019,     0.01019,
  0.01019,    0.01019,     0.01019,     0.01019,
  0.009984,   0.009984,    0.009984,    0.009984,
  0.009499,   0.009499,    0.009499,    0.009499,
  0.009162,   0.009162,    0.009162,    0.009162,
  0.008686,   0.008686,    0.008686,    0.008686,
  0.008066,   0.008066,    0.008066,    0.008066,
  0.007295,   0.007295,    0.007295,    0.007295,
  0.007057,   0.007057,    0.007057,    0.007057,
  0.007186,   0.007186,    0.007186,    0.007186,
  0.007033,   0.007033,    0.007033,    0.007033,
  0.006959,   0.006959,    0.006959,    0.006959,
  0.006759,   0.006759,    0.006759,    0.006759,
  0.006498,   0.006498,    0.006498,    0.006498,
  0.006301,   0.006301,    0.006301,    0.006301,
  0.006377,   0.006377,    0.006377,    0.006377,
  0.006629,   0.006629,    0.006629,    0.006629,
  0.00701,    0.00701,     0.00701,     0.00701,
  0.008136,   0.008136,    0.008136,    0.008136,
  0.009197,   0.009197,    0.009197,    0.009197,
  0.009446,   0.009446,    0.009446,    0.009446,
  0.009479,   0.009479,    0.009479,    0.009479,
  0.009519,   0.009519,    0.009519,    0.009519,
  0.009655,   0.009655,    0.009655,    0.009655,
  0.009843,   0.009843,    0.009843,    0.009843,
  0.009991,   0.009991,    0.009991,    0.009991,
  0.01008,    0.01008,     0.01008,     0.01008,
  0.009913,   0.009913,    0.009913,    0.009913,
  0.009653,   0.009653,    0.009653,    0.009653,
  0.009578,   0.009578,    0.009578,    0.009578,
  0.009647,   0.009647,    0.009647,    0.009647,
  0.009772,   0.009772,    0.009772,    0.009772,
  0.009759,   0.009759,    0.009759,    0.009759,
  0.009785,   0.009785,    0.009785,    0.009785,
  0.009905,   0.009905,    0.009905,    0.009905,
  0.009939,   0.009939,    0.009939,    0.009939,
  0.01,       0.01,        0.01,        0.01,
  0.01001,    0.01001,     0.01001,     0.01001,
  0.009933,   0.009933,    0.009933,    0.009933,
  0.009971,   0.009971,    0.009971,    0.009971,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.009984,   0.009984,    0.009984,    0.009984,
  0.01011,    0.01011,     0.01011,     0.01011,
  0.01021,    0.01021,     0.01021,     0.01021,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01059,    0.01059,     0.01059,     0.01059,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.009623,   0.009623,    0.009623,    0.009623,
  0.008753,   0.008753,    0.008753,    0.008753,
  0.007765,   0.007765,    0.007765,    0.007765,
  0.006692,   0.006692,    0.006692,    0.006692,
  0.005661,   0.005661,    0.005661,    0.005661,
  0.004962,   0.004962,    0.004962,    0.004962,
  0.004457,   0.004457,    0.004457,    0.004457,
  0.004269,   0.004269,    0.004269,    0.004269,
  0.004102,   0.004102,    0.004102,    0.004102,
  0.003363,   0.003363,    0.003363,    0.003363,
  0.003125,   0.003125,    0.003125,    0.003125,
  0.003372,   0.003372,    0.003372,    0.003372,
  0.003278,   0.003278,    0.003278,    0.003278,
  0.003131,   0.003131,    0.003131,    0.003131,
  0.003465,   0.003465,    0.003465,    0.003465,
  0.0039,     0.0039,      0.0039,      0.0039,
  0.003745,   0.003745,    0.003745,    0.003745,
  0.003533,   0.003533,    0.003533,    0.003533,
  0.003827,   0.003827,    0.003827,    0.003827,
  0.00451,    0.00451,     0.00451,     0.00451,
  0.005043,   0.005043,    0.005043,    0.005043,
  0.005338,   0.005338,    0.005338,    0.005338,
  0.00565,    0.00565,     0.00565,     0.00565,
  0.006088,   0.006088,    0.006088,    0.006088,
  0.00661,    0.00661,     0.00661,     0.00661,
  0.007052,   0.007052,    0.007052,    0.007052,
  0.007485,   0.007485,    0.007485,    0.007485,
  0.007803,   0.007803,    0.007803,    0.007803,
  0.007896,   0.007896,    0.007896,    0.007896,
  0.00793,    0.00793,     0.00793,     0.00793,
  0.007881,   0.007881,    0.007881,    0.007881,
  0.007711,   0.007711,    0.007711,    0.007711,
  0.007546,   0.007546,    0.007546,    0.007546,
  0.007384,   0.007384,    0.007384,    0.007384,
  0.00716,    0.00716,     0.00716,     0.00716,
  0.00697,    0.00697,     0.00697,     0.00697,
  0.006908,   0.006908,    0.006908,    0.006908,
  0.006881,   0.006881,    0.006881,    0.006881,
  0.006829,   0.006829,    0.006829,    0.006829,
  0.00682,    0.00682,     0.00682,     0.00682,
  0.006742,   0.006742,    0.006742,    0.006742,
  0.006594,   0.006594,    0.006594,    0.006594,
  0.00661,    0.00661,     0.00661,     0.00661,
  0.00679,    0.00679,     0.00679,     0.00679,
  0.007003,   0.007003,    0.007003,    0.007003,
  0.007201,   0.007201,    0.007201,    0.007201,
  0.007205,   0.007205,    0.007205,    0.007205,
  0.007004,   0.007004,    0.007004,    0.007004,
  0.006583,   0.006583,    0.006583,    0.006583,
  0.00581,    0.00581,     0.00581,     0.00581,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005771,   0.005771,    0.005771,    0.005771,
  0.005421,   0.005421,    0.005421,    0.005421,
  0.00503,    0.00503,     0.00503,     0.00503,
  0.005099,   0.005099,    0.005099,    0.005099,
  0.005282,   0.005282,    0.005282,    0.005282,
  0.004994,   0.004994,    0.004994,    0.004994,
  0.004619,   0.004619,    0.004619,    0.004619,
  0.004727,   0.004727,    0.004727,    0.004727,
  0.005191,   0.005191,    0.005191,    0.005191,
  0.005642,   0.005642,    0.005642,    0.005642,
  0.005792,   0.005792,    0.005792,    0.005792,
  0.005836,   0.005836,    0.005836,    0.005836,
  0.005945,   0.005945,    0.005945,    0.005945,
  0.006128,   0.006128,    0.006128,    0.006128,
  0.006429,   0.006429,    0.006429,    0.006429,
  0.006366,   0.006366,    0.006366,    0.006366,
  0.006084,   0.006084,    0.006084,    0.006084,
  0.006661,   0.006661,    0.006661,    0.006661,
  0.007351,   0.007351,    0.007351,    0.007351,
  0.007574,   0.007574,    0.007574,    0.007574,
  0.007855,   0.007855,    0.007855,    0.007855,
  0.008148,   0.008148,    0.008148,    0.008148,
  0.008453,   0.008453,    0.008453,    0.008453,
  0.008737,   0.008737,    0.008737,    0.008737,
  0.008997,   0.008997,    0.008997,    0.008997,
  0.009196,   0.009196,    0.009196,    0.009196,
  0.009276,   0.009276,    0.009276,    0.009276,
  0.009297,   0.009297,    0.009297,    0.009297,
  0.009319,   0.009319,    0.009319,    0.009319,
  0.009286,   0.009286,    0.009286,    0.009286,
  0.00927,    0.00927,     0.00927,     0.00927,
  0.009275,   0.009275,    0.009275,    0.009275,
  0.009263,   0.009263,    0.009263,    0.009263,
  0.009267,   0.009267,    0.009267,    0.009267,
  0.009267,   0.009267,    0.009267,    0.009267,
  0.00929,    0.00929,     0.00929,     0.00929,
  0.009357,   0.009357,    0.009357,    0.009357,
  0.009439,   0.009439,    0.009439,    0.009439,
  0.009443,   0.009443,    0.009443,    0.009443,
  0.009419,   0.009419,    0.009419,    0.009419,
  0.009471,   0.009471,    0.009471,    0.009471,
  0.009621,   0.009621,    0.009621,    0.009621,
  0.009825,   0.009825,    0.009825,    0.009825,
  0.009877,   0.009877,    0.009877,    0.009877,
  0.009669,   0.009669,    0.009669,    0.009669,
  0.009422,   0.009422,    0.009422,    0.009422,
  0.009177,   0.009177,    0.009177,    0.009177,
  0.00909,    0.00909,     0.00909,     0.00909,
  0.009232,   0.009232,    0.009232,    0.009232,
  0.009271,   0.009271,    0.009271,    0.009271,
  0.009243,   0.009243,    0.009243,    0.009243,
  0.009254,   0.009254,    0.009254,    0.009254,
  0.009254,   0.009254,    0.009254,    0.009254,
  0.009187,   0.009187,    0.009187,    0.009187,
  0.009097,   0.009097,    0.009097,    0.009097,
  0.008877,   0.008877,    0.008877,    0.008877,
  0.008619,   0.008619,    0.008619,    0.008619,
  0.008591,   0.008591,    0.008591,    0.008591,
  0.008577,   0.008577,    0.008577,    0.008577,
  0.008312,   0.008312,    0.008312,    0.008312,
  0.008079,   0.008079,    0.008079,    0.008079,
  0.008136,   0.008136,    0.008136,    0.008136,
  0.008245,   0.008245,    0.008245,    0.008245,
  0.008315,   0.008315,    0.008315,    0.008315,
  0.008407,   0.008407,    0.008407,    0.008407,
  0.008519,   0.008519,    0.008519,    0.008519,
  0.008656,   0.008656,    0.008656,    0.008656,
  0.009074,   0.009074,    0.009074,    0.009074,
  0.00955,    0.00955,     0.00955,     0.00955,
  0.009735,   0.009735,    0.009735,    0.009735,
  0.009881,   0.009881,    0.009881,    0.009881,
  0.01001,    0.01001,     0.01001,     0.01001,
  0.01005,    0.01005,     0.01005,     0.01005,
  0.01,       0.01,        0.01,        0.01,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.01012,    0.01012,     0.01012,     0.01012,
  0.01015,    0.01015,     0.01015,     0.01015,
  0.01,       0.01,        0.01,        0.01,
  0.009887,   0.009887,    0.009887,    0.009887,
  0.01004,    0.01004,     0.01004,     0.01004,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.009977,   0.009977,    0.009977,    0.009977,
  0.009839,   0.009839,    0.009839,    0.009839,
  0.009816,   0.009816,    0.009816,    0.009816,
  0.009879,   0.009879,    0.009879,    0.009879,
  0.00983,    0.00983,     0.00983,     0.00983,
  0.009867,   0.009867,    0.009867,    0.009867,
  0.009947,   0.009947,    0.009947,    0.009947,
  0.009994,   0.009994,    0.009994,    0.009994,
  0.01011,    0.01011,     0.01011,     0.01011,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.01041,    0.01041,     0.01041,     0.01041,
  0.01068,    0.01068,     0.01068,     0.01068,
  0.01103,    0.01103,     0.01103,     0.01103,
  0.0112,     0.0112,      0.0112,      0.0112,
  0.01113,    0.01113,     0.01113,     0.01113,
  0.01086,    0.01086,     0.01086,     0.01086,
  0.01066,    0.01066,     0.01066,     0.01066,
  0.01046,    0.01046,     0.01046,     0.01046,
  0.009945,   0.009945,    0.009945,    0.009945,
  0.009439,   0.009439,    0.009439,    0.009439,
  0.009057,   0.009057,    0.009057,    0.009057,
  0.008736,   0.008736,    0.008736,    0.008736,
  0.008538,   0.008538,    0.008538,    0.008538,
  0.008049,   0.008049,    0.008049,    0.008049,
  0.007468,   0.007468,    0.007468,    0.007468,
  0.007373,   0.007373,    0.007373,    0.007373,
  0.007468,   0.007468,    0.007468,    0.007468,
  0.007453,   0.007453,    0.007453,    0.007453,
  0.007342,   0.007342,    0.007342,    0.007342,
  0.007136,   0.007136,    0.007136,    0.007136,
  0.006994,   0.006994,    0.006994,    0.006994,
  0.007089,   0.007089,    0.007089,    0.007089,
  0.007415,   0.007415,    0.007415,    0.007415,
  0.007608,   0.007608,    0.007608,    0.007608,
  0.007715,   0.007715,    0.007715,    0.007715,
  0.007871,   0.007871,    0.007871,    0.007871,
  0.008299,   0.008299,    0.008299,    0.008299,
  0.008662,   0.008662,    0.008662,    0.008662,
  0.008718,   0.008718,    0.008718,    0.008718,
  0.008933,   0.008933,    0.008933,    0.008933,
  0.009076,   0.009076,    0.009076,    0.009076,
  0.009126,   0.009126,    0.009126,    0.009126,
  0.009126,   0.009126,    0.009126,    0.009126,
  0.009094,   0.009094,    0.009094,    0.009094,
  0.009079,   0.009079,    0.009079,    0.009079,
  0.009032,   0.009032,    0.009032,    0.009032,
  0.00905,    0.00905,     0.00905,     0.00905,
  0.009078,   0.009078,    0.009078,    0.009078,
  0.008993,   0.008993,    0.008993,    0.008993,
  0.009028,   0.009028,    0.009028,    0.009028,
  0.00956,    0.00956,     0.00956,     0.00956,
  0.01039,    0.01039,     0.01039,     0.01039,
  0.01109,    0.01109,     0.01109,     0.01109,
  0.01146,    0.01146,     0.01146,     0.01146,
  0.01152,    0.01152,     0.01152,     0.01152,
  0.01155,    0.01155,     0.01155,     0.01155,
  0.01165,    0.01165,     0.01165,     0.01165,
  0.01177,    0.01177,     0.01177,     0.01177,
  0.01185,    0.01185,     0.01185,     0.01185,
  0.01193,    0.01193,     0.01193,     0.01193,
  0.01206,    0.01206,     0.01206,     0.01206,
  0.01214,    0.01214,     0.01214,     0.01214,
  0.01212,    0.01212,     0.01212,     0.01212,
  0.01213,    0.01213,     0.01213,     0.01213,
  0.0119,     0.0119,      0.0119,      0.0119,
  0.0117,     0.0117,      0.0117,      0.0117,
  0.01186,    0.01186,     0.01186,     0.01186,
  0.01196,    0.01196,     0.01196,     0.01196,
  0.01193,    0.01193,     0.01193,     0.01193,
  0.01186,    0.01186,     0.01186,     0.01186,
  0.01183,    0.01183,     0.01183,     0.01183,
  0.01183,    0.01183,     0.01183,     0.01183,
  0.01183,    0.01183,     0.01183,     0.01183,
  0.0119,     0.0119,      0.0119,      0.0119,
  0.01203,    0.01203,     0.01203,     0.01203,
  0.01213,    0.01213,     0.01213,     0.01213,
  0.01219,    0.01219,     0.01219,     0.01219,
  0.01226,    0.01226,     0.01226,     0.01226,
  0.01233,    0.01233,     0.01233,     0.01233,
  0.01236,    0.01236,     0.01236,     0.01236,
  0.01236,    0.01236,     0.01236,     0.01236,
  0.01236,    0.01236,     0.01236,     0.01236,
  0.01233,    0.01233,     0.01233,     0.01233,
  0.01226,    0.01226,     0.01226,     0.01226,
  0.01219,    0.01219,     0.01219,     0.01219,
  0.01216,    0.01216,     0.01216,     0.01216,
  0.01213,    0.01213,     0.01213,     0.01213,
  0.01206,    0.01206,     0.01206,     0.01206,
  0.01203,    0.01203,     0.01203,     0.01203,
  0.01203,    0.01203,     0.01203,     0.01203,
  0.01203,    0.01203,     0.01203,     0.01203,
  0.01203,    0.01203,     0.01203,     0.01203,
  0.01199,    0.01199,     0.01199,     0.01199,
  0.01193,    0.01193,     0.01193,     0.01193,
  0.01186,    0.01186,     0.01186,     0.01186,
  0.01183,    0.01183,     0.01183,     0.01183,
  0.0118,     0.0118,      0.0118,      0.0118,
  0.01176,    0.01176,     0.01176,     0.01176,
  0.01176,    0.01176,     0.01176,     0.01176,
  0.01176,    0.01176,     0.01176,     0.01176,
  0.01176,    0.01176,     0.01176,     0.01176,
  0.01173,    0.01173,     0.01173,     0.01173,
  0.0117,     0.0117,      0.0117,      0.0117,
  0.01167,    0.01167,     0.01167,     0.01167,
  0.01164,    0.01164,     0.01164,     0.01164,
  0.0116,     0.0116,      0.0116,      0.0116,
  0.01154,    0.01154,     0.01154,     0.01154,
  0.0116,     0.0116,      0.0116,      0.0116,
  0.0118,     0.0118,      0.0118,      0.0118,
  0.01199,    0.01199,     0.01199,     0.01199,
  0.0123,     0.0123,      0.0123,      0.0123,
  0.01264,    0.01264,     0.01264,     0.01264,
  0.01299,    0.01299,     0.01299,     0.01299,
  0.01342,    0.01342,     0.01342,     0.01342,
  0.01348,    0.01348,     0.01348,     0.01348,
  0.01322,    0.01322,     0.01322,     0.01322,
  0.01294,    0.01294,     0.01294,     0.01294,
  0.01272,    0.01272,     0.01272,     0.01272,
  0.01267,    0.01267,     0.01267,     0.01267,
  0.01255,    0.01255,     0.01255,     0.01255,
  0.01237,    0.01237,     0.01237,     0.01237,
  0.01212,    0.01212,     0.01212,     0.01212,
  0.01198,    0.01198,     0.01198,     0.01198,
  0.01206,    0.01206,     0.01206,     0.01206,
  0.01215,    0.01215,     0.01215,     0.01215,
  0.01236,    0.01236,     0.01236,     0.01236,
  0.01262,    0.01262,     0.01262,     0.01262,
  0.01284,    0.01284,     0.01284,     0.01284,
  0.01295,    0.01295,     0.01295,     0.01295,
  0.01301,    0.01301,     0.01301,     0.01301,
  0.01322,    0.01322,     0.01322,     0.01322,
  0.01331,    0.01331,     0.01331,     0.01331,
  0.01316,    0.01316,     0.01316,     0.01316,
  0.01297,    0.01297,     0.01297,     0.01297,
  0.01284,    0.01284,     0.01284,     0.01284,
  0.01272,    0.01272,     0.01272,     0.01272,
  0.01261,    0.01261,     0.01261,     0.01261,
  0.01261,    0.01261,     0.01261,     0.01261,
  0.01263,    0.01263,     0.01263,     0.01263,
  0.01262,    0.01262,     0.01262,     0.01262,
  0.01259,    0.01259,     0.01259,     0.01259,
  0.01255,    0.01255,     0.01255,     0.01255,
  0.01254,    0.01254,     0.01254,     0.01254,
  0.01249,    0.01249,     0.01249,     0.01249,
  0.01244,    0.01244,     0.01244,     0.01244,
  0.01243,    0.01243,     0.01243,     0.01243,
  0.01242,    0.01242,     0.01242,     0.01242,
  0.01233,    0.01233,     0.01233,     0.01233,
  0.01222,    0.01222,     0.01222,     0.01222,
  0.01215,    0.01215,     0.01215,     0.01215,
  0.01207,    0.01207,     0.01207,     0.01207,
  0.01208,    0.01208,     0.01208,     0.01208,
  0.01216,    0.01216,     0.01216,     0.01216,
  0.01217,    0.01217,     0.01217,     0.01217,
  0.01211,    0.01211,     0.01211,     0.01211,
  0.0121,     0.0121,      0.0121,      0.0121,
  0.01221,    0.01221,     0.01221,     0.01221,
  0.01244,    0.01244,     0.01244,     0.01244,
  0.01256,    0.01256,     0.01256,     0.01256,
  0.01223,    0.01223,     0.01223,     0.01223,
  0.01178,    0.01178,     0.01178,     0.01178,
  0.01165,    0.01165,     0.01165,     0.01165,
  0.01166,    0.01166,     0.01166,     0.01166,
  0.01142,    0.01142,     0.01142,     0.01142,
  0.01107,    0.01107,     0.01107,     0.01107,
  0.0109,     0.0109,      0.0109,      0.0109,
  0.01086,    0.01086,     0.01086,     0.01086,
  0.01099,    0.01099,     0.01099,     0.01099,
  0.01098,    0.01098,     0.01098,     0.01098,
  0.01084,    0.01084,     0.01084,     0.01084,
  0.01079,    0.01079,     0.01079,     0.01079,
  0.01077,    0.01077,     0.01077,     0.01077,
  0.01067,    0.01067,     0.01067,     0.01067,
  0.0106,     0.0106,      0.0106,      0.0106,
  0.01073,    0.01073,     0.01073,     0.01073,
  0.01093,    0.01093,     0.01093,     0.01093,
  0.0111,     0.0111,      0.0111,      0.0111,
  0.01109,    0.01109,     0.01109,     0.01109,
  0.01124,    0.01124,     0.01124,     0.01124,
  0.01168,    0.01168,     0.01168,     0.01168,
  0.01206,    0.01206,     0.01206,     0.01206,
  0.01221,    0.01221,     0.01221,     0.01221,
  0.01231,    0.01231,     0.01231,     0.01231,
  0.01255,    0.01255,     0.01255,     0.01255,
  0.0127,     0.0127,      0.0127,      0.0127,
  0.01273,    0.01273,     0.01273,     0.01273,
  0.01263,    0.01263,     0.01263,     0.01263,
  0.0123,     0.0123,      0.0123,      0.0123,
  0.01205,    0.01205,     0.01205,     0.01205,
  0.01199,    0.01199,     0.01199,     0.01199,
  0.01203,    0.01203,     0.01203,     0.01203,
  0.01216,    0.01216,     0.01216,     0.01216,
  0.01226,    0.01226,     0.01226,     0.01226,
  0.0123,     0.0123,      0.0123,      0.0123,
  0.01226,    0.01226,     0.01226,     0.01226,
  0.01213,    0.01213,     0.01213,     0.01213,
  0.01196,    0.01196,     0.01196,     0.01196,
  0.01186,    0.01186,     0.01186,     0.01186,
  0.01183,    0.01183,     0.01183,     0.01183,
  0.0119,     0.0119,      0.0119,      0.0119,
  0.01206,    0.01206,     0.01206,     0.01206,
  0.01233,    0.01233,     0.01233,     0.01233,
  0.01271,    0.01271,     0.01271,     0.01271,
  0.01317,    0.01317,     0.01317,     0.01317,
  0.01339,    0.01339,     0.01339,     0.01339,
  0.01342,    0.01342,     0.01342,     0.01342,
  0.01339,    0.01339,     0.01339,     0.01339,
  0.01312,    0.01312,     0.01312,     0.01312,
  0.01293,    0.01293,     0.01293,     0.01293,
  0.01272,    0.01272,     0.01272,     0.01272,
  0.01192,    0.01192,     0.01192,     0.01192,
  0.01145,    0.01145,     0.01145,     0.01145,
  0.01133,    0.01133,     0.01133,     0.01133,
  0.01057,    0.01057,     0.01057,     0.01057,
  0.009671,   0.009671,    0.009671,    0.009671,
  0.009204,   0.009204,    0.009204,    0.009204,
  0.009282,   0.009282,    0.009282,    0.009282,
  0.009796,   0.009796,    0.009796,    0.009796,
  0.01038,    0.01038,     0.01038,     0.01038,
  0.01107,    0.01107,     0.01107,     0.01107,
  0.01174,    0.01174,     0.01174,     0.01174,
  0.012,      0.012,       0.012,       0.012,
  0.01203,    0.01203,     0.01203,     0.01203,
  0.01209,    0.01209,     0.01209,     0.01209,
  0.01216,    0.01216,     0.01216,     0.01216,
  0.01216,    0.01216,     0.01216,     0.01216,
  0.01216,    0.01216,     0.01216,     0.01216,
  0.01216,    0.01216,     0.01216,     0.01216,
  0.01213,    0.01213,     0.01213,     0.01213,
  0.01206,    0.01206,     0.01206,     0.01206,
  0.01203,    0.01203,     0.01203,     0.01203,
  0.0119,     0.0119,      0.0119,      0.0119,
  0.01167,    0.01167,     0.01167,     0.01167,
  0.01148,    0.01148,     0.01148,     0.01148,
  0.01132,    0.01132,     0.01132,     0.01132,
  0.01125,    0.01125,     0.01125,     0.01125,
  0.01125,    0.01125,     0.01125,     0.01125,
  0.01122,    0.01122,     0.01122,     0.01122,
  0.01119,    0.01119,     0.01119,     0.01119,
  0.01116,    0.01116,     0.01116,     0.01116,
  0.01107,    0.01107,     0.01107,     0.01107,
  0.01098,    0.01098,     0.01098,     0.01098,
  0.01094,    0.01094,     0.01094,     0.01094,
  0.01101,    0.01101,     0.01101,     0.01101,
  0.0111,     0.0111,      0.0111,      0.0111,
  0.01116,    0.01116,     0.01116,     0.01116,
  0.01119,    0.01119,     0.01119,     0.01119,
  0.01119,    0.01119,     0.01119,     0.01119,
  0.01119,    0.01119,     0.01119,     0.01119,
  0.01119,    0.01119,     0.01119,     0.01119,
  0.01125,    0.01125,     0.01125,     0.01125,
  0.01141,    0.01141,     0.01141,     0.01141,
  0.0116,     0.0116,      0.0116,      0.0116,
  0.0118,     0.0118,      0.0118,      0.0118,
  0.01187,    0.01187,     0.01187,     0.01187,
  0.01172,    0.01172,     0.01172,     0.01172,
  0.01161,    0.01161,     0.01161,     0.01161,
  0.01147,    0.01147,     0.01147,     0.01147,
  0.01129,    0.01129,     0.01129,     0.01129,
  0.01131,    0.01131,     0.01131,     0.01131,
  0.01096,    0.01096,     0.01096,     0.01096,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.01092,    0.01092,     0.01092,     0.01092,
  0.0111,     0.0111,      0.0111,      0.0111,
  0.01094,    0.01094,     0.01094,     0.01094,
  0.0108,     0.0108,      0.0108,      0.0108,
  0.01088,    0.01088,     0.01088,     0.01088,
  0.0109,     0.0109,      0.0109,      0.0109,
  0.01086,    0.01086,     0.01086,     0.01086,
  0.01089,    0.01089,     0.01089,     0.01089,
  0.0108,     0.0108,      0.0108,      0.0108,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01047,    0.01047,     0.01047,     0.01047,
  0.01086,    0.01086,     0.01086,     0.01086,
  0.01107,    0.01107,     0.01107,     0.01107,
  0.01094,    0.01094,     0.01094,     0.01094,
  0.01082,    0.01082,     0.01082,     0.01082,
  0.01079,    0.01079,     0.01079,     0.01079,
  0.01067,    0.01067,     0.01067,     0.01067,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01047,    0.01047,     0.01047,     0.01047,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.009758,   0.009758,    0.009758,    0.009758,
  0.009481,   0.009481,    0.009481,    0.009481,
  0.009563,   0.009563,    0.009563,    0.009563,
  0.009617,   0.009617,    0.009617,    0.009617,
  0.009644,   0.009644,    0.009644,    0.009644,
  0.009644,   0.009644,    0.009644,    0.009644,
  0.009617,   0.009617,    0.009617,    0.009617,
  0.009644,   0.009644,    0.009644,    0.009644,
  0.009563,   0.009563,    0.009563,    0.009563,
  0.009401,   0.009401,    0.009401,    0.009401,
  0.009401,   0.009401,    0.009401,    0.009401,
  0.009563,   0.009563,    0.009563,    0.009563,
  0.009754,   0.009754,    0.009754,    0.009754,
  0.009893,   0.009893,    0.009893,    0.009893,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.01023,    0.01023,     0.01023,     0.01023,
  0.01041,    0.01041,     0.01041,     0.01041,
  0.01067,    0.01067,     0.01067,     0.01067,
  0.01085,    0.01085,     0.01085,     0.01085,
  0.01116,    0.01116,     0.01116,     0.01116,
  0.01125,    0.01125,     0.01125,     0.01125,
  0.0109,     0.0109,      0.0109,      0.0109,
  0.01062,    0.01062,     0.01062,     0.01062,
  0.01053,    0.01053,     0.01053,     0.01053,
  0.01038,    0.01038,     0.01038,     0.01038,
  0.01002,    0.01002,     0.01002,     0.01002,
  0.009637,   0.009637,    0.009637,    0.009637,
  0.009304,   0.009304,    0.009304,    0.009304,
  0.009288,   0.009288,    0.009288,    0.009288,
  0.009191,   0.009191,    0.009191,    0.009191,
  0.009078,   0.009078,    0.009078,    0.009078,
  0.009475,   0.009475,    0.009475,    0.009475,
  0.009932,   0.009932,    0.009932,    0.009932,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01072,    0.01072,     0.01072,     0.01072,
  0.011,      0.011,       0.011,       0.011,
  0.01122,    0.01122,     0.01122,     0.01122,
  0.01125,    0.01125,     0.01125,     0.01125,
  0.01107,    0.01107,     0.01107,     0.01107,
  0.01091,    0.01091,     0.01091,     0.01091,
  0.01082,    0.01082,     0.01082,     0.01082,
  0.0107,     0.0107,      0.0107,      0.0107,
  0.01067,    0.01067,     0.01067,     0.01067,
  0.01073,    0.01073,     0.01073,     0.01073,
  0.01082,    0.01082,     0.01082,     0.01082,
  0.01091,    0.01091,     0.01091,     0.01091,
  0.01091,    0.01091,     0.01091,     0.01091,
  0.01085,    0.01085,     0.01085,     0.01085,
  0.01081,    0.01081,     0.01081,     0.01081,
  0.01082,    0.01082,     0.01082,     0.01082,
  0.01082,    0.01082,     0.01082,     0.01082,
  0.01082,    0.01082,     0.01082,     0.01082,
  0.01079,    0.01079,     0.01079,     0.01079,
  0.0107,     0.0107,      0.0107,      0.0107,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.0105,     0.0105,      0.0105,      0.0105,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01041,    0.01041,     0.01041,     0.01041,
  0.01035,    0.01035,     0.01035,     0.01035,
  0.01029,    0.01029,     0.01029,     0.01029,
  0.01029,    0.01029,     0.01029,     0.01029,
  0.01029,    0.01029,     0.01029,     0.01029,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01038,    0.01038,     0.01038,     0.01038,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01035,    0.01035,     0.01035,     0.01035,
  0.01015,    0.01015,     0.01015,     0.01015,
  0.01012,    0.01012,     0.01012,     0.01012,
  0.01026,    0.01026,     0.01026,     0.01026,
  0.01027,    0.01027,     0.01027,     0.01027,
  0.0102,     0.0102,      0.0102,      0.0102,
  0.01017,    0.01017,     0.01017,     0.01017,
  0.009982,   0.009982,    0.009982,    0.009982,
  0.009547,   0.009547,    0.009547,    0.009547,
  0.009041,   0.009041,    0.009041,    0.009041,
  0.008846,   0.008846,    0.008846,    0.008846,
  0.009098,   0.009098,    0.009098,    0.009098,
  0.009374,   0.009374,    0.009374,    0.009374,
  0.00943,    0.00943,     0.00943,     0.00943,
  0.009402,   0.009402,    0.009402,    0.009402,
  0.009442,   0.009442,    0.009442,    0.009442,
  0.009448,   0.009448,    0.009448,    0.009448,
  0.008631,   0.008631,    0.008631,    0.008631,
  0.007734,   0.007734,    0.007734,    0.007734,
  0.007687,   0.007687,    0.007687,    0.007687,
  0.00784,    0.00784,     0.00784,     0.00784,
  0.00804,    0.00804,     0.00804,     0.00804,
  0.008281,   0.008281,    0.008281,    0.008281,
  0.008418,   0.008418,    0.008418,    0.008418,
  0.008513,   0.008513,    0.008513,    0.008513,
  0.008571,   0.008571,    0.008571,    0.008571,
  0.008541,   0.008541,    0.008541,    0.008541,
  0.00842,    0.00842,     0.00842,     0.00842,
  0.008105,   0.008105,    0.008105,    0.008105,
  0.007858,   0.007858,    0.007858,    0.007858,
  0.007877,   0.007877,    0.007877,    0.007877,
  0.00795,    0.00795,     0.00795,     0.00795,
  0.008003,   0.008003,    0.008003,    0.008003,
  0.008056,   0.008056,    0.008056,    0.008056,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008139,   0.008139,    0.008139,    0.008139,
  0.008265,   0.008265,    0.008265,    0.008265,
  0.008397,   0.008397,    0.008397,    0.008397,
  0.008391,   0.008391,    0.008391,    0.008391,
  0.00835,    0.00835,     0.00835,     0.00835,
  0.00825,    0.00825,     0.00825,     0.00825,
  0.008177,   0.008177,    0.008177,    0.008177,
  0.00819,    0.00819,     0.00819,     0.00819,
  0.008192,   0.008192,    0.008192,    0.008192,
  0.008196,   0.008196,    0.008196,    0.008196,
  0.00815,    0.00815,     0.00815,     0.00815,
  0.008137,   0.008137,    0.008137,    0.008137,
  0.008089,   0.008089,    0.008089,    0.008089,
  0.008071,   0.008071,    0.008071,    0.008071,
  0.008059,   0.008059,    0.008059,    0.008059,
  0.007925,   0.007925,    0.007925,    0.007925,
  0.007856,   0.007856,    0.007856,    0.007856,
  0.007953,   0.007953,    0.007953,    0.007953,
  0.008414,   0.008414,    0.008414,    0.008414,
  0.008414,   0.008414,    0.008414,    0.008414,
  0.008027,   0.008027,    0.008027,    0.008027,
  0.0079,     0.0079,      0.0079,      0.0079,
  0.007808,   0.007808,    0.007808,    0.007808,
  0.007796,   0.007796,    0.007796,    0.007796,
  0.007435,   0.007435,    0.007435,    0.007435,
  0.007166,   0.007166,    0.007166,    0.007166,
  0.007398,   0.007398,    0.007398,    0.007398,
  0.007825,   0.007825,    0.007825,    0.007825,
  0.008226,   0.008226,    0.008226,    0.008226,
  0.008358,   0.008358,    0.008358,    0.008358,
  0.008454,   0.008454,    0.008454,    0.008454,
  0.008562,   0.008562,    0.008562,    0.008562,
  0.00852,    0.00852,     0.00852,     0.00852,
  0.008495,   0.008495,    0.008495,    0.008495,
  0.008371,   0.008371,    0.008371,    0.008371,
  0.008195,   0.008195,    0.008195,    0.008195,
  0.00809,    0.00809,     0.00809,     0.00809,
  0.007972,   0.007972,    0.007972,    0.007972,
  0.007886,   0.007886,    0.007886,    0.007886,
  0.007783,   0.007783,    0.007783,    0.007783,
  0.007634,   0.007634,    0.007634,    0.007634,
  0.007518,   0.007518,    0.007518,    0.007518,
  0.007475,   0.007475,    0.007475,    0.007475,
  0.007378,   0.007378,    0.007378,    0.007378,
  0.007262,   0.007262,    0.007262,    0.007262,
  0.007208,   0.007208,    0.007208,    0.007208,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007155,   0.007155,    0.007155,    0.007155,
  0.007209,   0.007209,    0.007209,    0.007209,
  0.007305,   0.007305,    0.007305,    0.007305,
  0.00738,    0.00738,     0.00738,     0.00738,
  0.007481,   0.007481,    0.007481,    0.007481,
  0.007633,   0.007633,    0.007633,    0.007633,
  0.00784,    0.00784,     0.00784,     0.00784,
  0.008087,   0.008087,    0.008087,    0.008087,
  0.008276,   0.008276,    0.008276,    0.008276,
  0.00844,    0.00844,     0.00844,     0.00844,
  0.008556,   0.008556,    0.008556,    0.008556,
  0.008552,   0.008552,    0.008552,    0.008552,
  0.008539,   0.008539,    0.008539,    0.008539,
  0.008641,   0.008641,    0.008641,    0.008641,
  0.008893,   0.008893,    0.008893,    0.008893,
  0.009228,   0.009228,    0.009228,    0.009228,
  0.009414,   0.009414,    0.009414,    0.009414,
  0.009311,   0.009311,    0.009311,    0.009311,
  0.009188,   0.009188,    0.009188,    0.009188,
  0.009182,   0.009182,    0.009182,    0.009182,
  0.009242,   0.009242,    0.009242,    0.009242,
  0.009466,   0.009466,    0.009466,    0.009466,
  0.009792,   0.009792,    0.009792,    0.009792,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.01021,    0.01021,     0.01021,     0.01021,
  0.0103,     0.0103,      0.0103,      0.0103,
  0.01038,    0.01038,     0.01038,     0.01038,
  0.01051,    0.01051,     0.01051,     0.01051,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.01058,    0.01058,     0.01058,     0.01058,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.01067,    0.01067,     0.01067,     0.01067,
  0.0107,     0.0107,      0.0107,      0.0107,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.01034,    0.01034,     0.01034,     0.01034,
  0.00995,    0.00995,     0.00995,     0.00995,
  0.009738,   0.009738,    0.009738,    0.009738,
  0.009549,   0.009549,    0.009549,    0.009549,
  0.009337,   0.009337,    0.009337,    0.009337,
  0.009281,   0.009281,    0.009281,    0.009281,
  0.009316,   0.009316,    0.009316,    0.009316,
  0.009291,   0.009291,    0.009291,    0.009291,
  0.009266,   0.009266,    0.009266,    0.009266,
  0.009274,   0.009274,    0.009274,    0.009274,
  0.009215,   0.009215,    0.009215,    0.009215,
  0.009179,   0.009179,    0.009179,    0.009179,
  0.009228,   0.009228,    0.009228,    0.009228,
  0.009232,   0.009232,    0.009232,    0.009232,
  0.00914,    0.00914,     0.00914,     0.00914,
  0.009091,   0.009091,    0.009091,    0.009091,
  0.008895,   0.008895,    0.008895,    0.008895,
  0.008577,   0.008577,    0.008577,    0.008577,
  0.008264,   0.008264,    0.008264,    0.008264,
  0.008143,   0.008143,    0.008143,    0.008143,
  0.008219,   0.008219,    0.008219,    0.008219,
  0.008196,   0.008196,    0.008196,    0.008196,
  0.008162,   0.008162,    0.008162,    0.008162,
  0.008175,   0.008175,    0.008175,    0.008175,
  0.008219,   0.008219,    0.008219,    0.008219,
  0.008172,   0.008172,    0.008172,    0.008172,
  0.008144,   0.008144,    0.008144,    0.008144,
  0.008089,   0.008089,    0.008089,    0.008089,
  0.008188,   0.008188,    0.008188,    0.008188,
  0.008491,   0.008491,    0.008491,    0.008491,
  0.008692,   0.008692,    0.008692,    0.008692,
  0.00878,    0.00878,     0.00878,     0.00878,
  0.008803,   0.008803,    0.008803,    0.008803,
  0.008831,   0.008831,    0.008831,    0.008831,
  0.008953,   0.008953,    0.008953,    0.008953,
  0.009078,   0.009078,    0.009078,    0.009078,
  0.009165,   0.009165,    0.009165,    0.009165,
  0.009322,   0.009322,    0.009322,    0.009322,
  0.00941,    0.00941,     0.00941,     0.00941,
  0.009279,   0.009279,    0.009279,    0.009279,
  0.009092,   0.009092,    0.009092,    0.009092,
  0.009024,   0.009024,    0.009024,    0.009024,
  0.009104,   0.009104,    0.009104,    0.009104,
  0.009251,   0.009251,    0.009251,    0.009251,
  0.009351,   0.009351,    0.009351,    0.009351,
  0.009485,   0.009485,    0.009485,    0.009485,
  0.009672,   0.009672,    0.009672,    0.009672,
  0.009823,   0.009823,    0.009823,    0.009823,
  0.009944,   0.009944,    0.009944,    0.009944,
  0.01007,    0.01007,     0.01007,     0.01007,
  0.01019,    0.01019,     0.01019,     0.01019,
  0.01028,    0.01028,     0.01028,     0.01028,
  0.01037,    0.01037,     0.01037,     0.01037,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.0105,     0.0105,      0.0105,      0.0105,
  0.01057,    0.01057,     0.01057,     0.01057,
  0.01057,    0.01057,     0.01057,     0.01057,
  0.01058,    0.01058,     0.01058,     0.01058,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.01038,    0.01038,     0.01038,     0.01038,
  0.009869,   0.009869,    0.009869,    0.009869,
  0.009497,   0.009497,    0.009497,    0.009497,
  0.009193,   0.009193,    0.009193,    0.009193,
  0.008616,   0.008616,    0.008616,    0.008616,
  0.00831,    0.00831,     0.00831,     0.00831,
  0.008586,   0.008586,    0.008586,    0.008586,
  0.008724,   0.008724,    0.008724,    0.008724,
  0.008619,   0.008619,    0.008619,    0.008619,
  0.008504,   0.008504,    0.008504,    0.008504,
  0.008245,   0.008245,    0.008245,    0.008245,
  0.007861,   0.007861,    0.007861,    0.007861,
  0.007609,   0.007609,    0.007609,    0.007609,
  0.007467,   0.007467,    0.007467,    0.007467,
  0.007347,   0.007347,    0.007347,    0.007347,
  0.007315,   0.007315,    0.007315,    0.007315,
  0.007288,   0.007288,    0.007288,    0.007288,
  0.00725,    0.00725,     0.00725,     0.00725,
  0.007436,   0.007436,    0.007436,    0.007436,
  0.007642,   0.007642,    0.007642,    0.007642,
  0.007718,   0.007718,    0.007718,    0.007718,
  0.007979,   0.007979,    0.007979,    0.007979,
  0.008307,   0.008307,    0.008307,    0.008307,
  0.00858,    0.00858,     0.00858,     0.00858,
  0.008989,   0.008989,    0.008989,    0.008989,
  0.009311,   0.009311,    0.009311,    0.009311,
  0.009583,   0.009583,    0.009583,    0.009583,
  0.009798,   0.009798,    0.009798,    0.009798,
  0.009816,   0.009816,    0.009816,    0.009816,
  0.00983,    0.00983,     0.00983,     0.00983,
  0.009809,   0.009809,    0.009809,    0.009809,
  0.009727,   0.009727,    0.009727,    0.009727,
  0.009617,   0.009617,    0.009617,    0.009617,
  0.009429,   0.009429,    0.009429,    0.009429,
  0.009164,   0.009164,    0.009164,    0.009164,
  0.008956,   0.008956,    0.008956,    0.008956,
  0.008854,   0.008854,    0.008854,    0.008854,
  0.008754,   0.008754,    0.008754,    0.008754,
  0.008531,   0.008531,    0.008531,    0.008531,
  0.008336,   0.008336,    0.008336,    0.008336,
  0.008216,   0.008216,    0.008216,    0.008216,
  0.008122,   0.008122,    0.008122,    0.008122,
  0.008122,   0.008122,    0.008122,    0.008122,
  0.008169,   0.008169,    0.008169,    0.008169,
  0.008216,   0.008216,    0.008216,    0.008216,
  0.008264,   0.008264,    0.008264,    0.008264,
  0.008312,   0.008312,    0.008312,    0.008312,
  0.008408,   0.008408,    0.008408,    0.008408,
  0.00853,    0.00853,     0.00853,     0.00853,
  0.008679,   0.008679,    0.008679,    0.008679,
  0.008829,   0.008829,    0.008829,    0.008829,
  0.009008,   0.009008,    0.009008,    0.009008,
  0.009184,   0.009184,    0.009184,    0.009184,
  0.009217,   0.009217,    0.009217,    0.009217,
  0.009275,   0.009275,    0.009275,    0.009275,
  0.009324,   0.009324,    0.009324,    0.009324,
  0.009214,   0.009214,    0.009214,    0.009214,
  0.008906,   0.008906,    0.008906,    0.008906,
  0.008457,   0.008457,    0.008457,    0.008457,
  0.008139,   0.008139,    0.008139,    0.008139,
  0.007901,   0.007901,    0.007901,    0.007901,
  0.007539,   0.007539,    0.007539,    0.007539,
  0.007334,   0.007334,    0.007334,    0.007334,
  0.007274,   0.007274,    0.007274,    0.007274,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007044,   0.007044,    0.007044,    0.007044,
  0.007318,   0.007318,    0.007318,    0.007318,
  0.007675,   0.007675,    0.007675,    0.007675,
  0.007937,   0.007937,    0.007937,    0.007937,
  0.008551,   0.008551,    0.008551,    0.008551,
  0.009176,   0.009176,    0.009176,    0.009176,
  0.009366,   0.009366,    0.009366,    0.009366,
  0.009375,   0.009375,    0.009375,    0.009375,
  0.009493,   0.009493,    0.009493,    0.009493,
  0.009521,   0.009521,    0.009521,    0.009521,
  0.009366,   0.009366,    0.009366,    0.009366,
  0.009275,   0.009275,    0.009275,    0.009275,
  0.009203,   0.009203,    0.009203,    0.009203,
  0.009127,   0.009127,    0.009127,    0.009127,
  0.009032,   0.009032,    0.009032,    0.009032,
  0.008907,   0.008907,    0.008907,    0.008907,
  0.008856,   0.008856,    0.008856,    0.008856,
  0.008711,   0.008711,    0.008711,    0.008711,
  0.008572,   0.008572,    0.008572,    0.008572,
  0.008482,   0.008482,    0.008482,    0.008482,
  0.008384,   0.008384,    0.008384,    0.008384,
  0.008265,   0.008265,    0.008265,    0.008265,
  0.008169,   0.008169,    0.008169,    0.008169,
  0.008169,   0.008169,    0.008169,    0.008169,
  0.008122,   0.008122,    0.008122,    0.008122,
  0.008052,   0.008052,    0.008052,    0.008052,
  0.008075,   0.008075,    0.008075,    0.008075,
  0.008052,   0.008052,    0.008052,    0.008052,
  0.007959,   0.007959,    0.007959,    0.007959,
  0.007913,   0.007913,    0.007913,    0.007913,
  0.008006,   0.008006,    0.008006,    0.008006,
  0.008313,   0.008313,    0.008313,    0.008313,
  0.008757,   0.008757,    0.008757,    0.008757,
  0.009317,   0.009317,    0.009317,    0.009317,
  0.009529,   0.009529,    0.009529,    0.009529,
  0.00938,    0.00938,     0.00938,     0.00938,
  0.009114,   0.009114,    0.009114,    0.009114,
  0.008685,   0.008685,    0.008685,    0.008685,
  0.008353,   0.008353,    0.008353,    0.008353,
  0.008208,   0.008208,    0.008208,    0.008208,
  0.007976,   0.007976,    0.007976,    0.007976,
  0.007551,   0.007551,    0.007551,    0.007551,
  0.00726,    0.00726,     0.00726,     0.00726,
  0.007169,   0.007169,    0.007169,    0.007169,
  0.007025,   0.007025,    0.007025,    0.007025,
  0.007007,   0.007007,    0.007007,    0.007007,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.007038,   0.007038,    0.007038,    0.007038,
  0.006932,   0.006932,    0.006932,    0.006932,
  0.006774,   0.006774,    0.006774,    0.006774,
  0.006961,   0.006961,    0.006961,    0.006961,
  0.007441,   0.007441,    0.007441,    0.007441,
  0.007757,   0.007757,    0.007757,    0.007757,
  0.007767,   0.007767,    0.007767,    0.007767,
  0.007784,   0.007784,    0.007784,    0.007784,
  0.008079,   0.008079,    0.008079,    0.008079,
  0.008423,   0.008423,    0.008423,    0.008423,
  0.008496,   0.008496,    0.008496,    0.008496,
  0.008478,   0.008478,    0.008478,    0.008478,
  0.00852,    0.00852,     0.00852,     0.00852,
  0.008524,   0.008524,    0.008524,    0.008524,
  0.008532,   0.008532,    0.008532,    0.008532,
  0.008538,   0.008538,    0.008538,    0.008538,
  0.008572,   0.008572,    0.008572,    0.008572,
  0.008641,   0.008641,    0.008641,    0.008641,
  0.008882,   0.008882,    0.008882,    0.008882,
  0.009109,   0.009109,    0.009109,    0.009109,
  0.00918,    0.00918,     0.00918,     0.00918,
  0.009212,   0.009212,    0.009212,    0.009212,
  0.009162,   0.009162,    0.009162,    0.009162,
  0.009157,   0.009157,    0.009157,    0.009157,
  0.009189,   0.009189,    0.009189,    0.009189,
  0.009117,   0.009117,    0.009117,    0.009117,
  0.009069,   0.009069,    0.009069,    0.009069,
  0.009176,   0.009176,    0.009176,    0.009176,
  0.009288,   0.009288,    0.009288,    0.009288,
  0.009319,   0.009319,    0.009319,    0.009319,
  0.009319,   0.009319,    0.009319,    0.009319,
  0.009432,   0.009432,    0.009432,    0.009432,
  0.009632,   0.009632,    0.009632,    0.009632,
  0.009853,   0.009853,    0.009853,    0.009853,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.01016,    0.01016,     0.01016,     0.01016,
  0.009998,   0.009998,    0.009998,    0.009998,
  0.009839,   0.009839,    0.009839,    0.009839,
  0.009684,   0.009684,    0.009684,    0.009684,
  0.009519,   0.009519,    0.009519,    0.009519,
  0.00926,    0.00926,     0.00926,     0.00926,
  0.008633,   0.008633,    0.008633,    0.008633,
  0.008323,   0.008323,    0.008323,    0.008323,
  0.008429,   0.008429,    0.008429,    0.008429,
  0.008022,   0.008022,    0.008022,    0.008022,
  0.007532,   0.007532,    0.007532,    0.007532,
  0.007501,   0.007501,    0.007501,    0.007501,
  0.007696,   0.007696,    0.007696,    0.007696,
  0.007854,   0.007854,    0.007854,    0.007854,
  0.007956,   0.007956,    0.007956,    0.007956,
  0.008194,   0.008194,    0.008194,    0.008194,
  0.008215,   0.008215,    0.008215,    0.008215,
  0.008238,   0.008238,    0.008238,    0.008238,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.007877,   0.007877,    0.007877,    0.007877,
  0.008141,   0.008141,    0.008141,    0.008141,
  0.008391,   0.008391,    0.008391,    0.008391,
  0.008496,   0.008496,    0.008496,    0.008496,
  0.008644,   0.008644,    0.008644,    0.008644,
  0.009019,   0.009019,    0.009019,    0.009019,
  0.009303,   0.009303,    0.009303,    0.009303,
  0.009343,   0.009343,    0.009343,    0.009343,
  0.00934,    0.00934,     0.00934,     0.00934,
  0.009363,   0.009363,    0.009363,    0.009363,
  0.009514,   0.009514,    0.009514,    0.009514,
  0.009666,   0.009666,    0.009666,    0.009666,
  0.009764,   0.009764,    0.009764,    0.009764,
  0.009804,   0.009804,    0.009804,    0.009804,
  0.00987,    0.00987,     0.00987,     0.00987,
  0.009904,   0.009904,    0.009904,    0.009904,
  0.009855,   0.009855,    0.009855,    0.009855,
  0.009806,   0.009806,    0.009806,    0.009806,
  0.009782,   0.009782,    0.009782,    0.009782,
  0.009699,   0.009699,    0.009699,    0.009699,
  0.009509,   0.009509,    0.009509,    0.009509,
  0.009321,   0.009321,    0.009321,    0.009321,
  0.009189,   0.009189,    0.009189,    0.009189,
  0.008983,   0.008983,    0.008983,    0.008983,
  0.008779,   0.008779,    0.008779,    0.008779,
  0.008829,   0.008829,    0.008829,    0.008829,
  0.009086,   0.009086,    0.009086,    0.009086,
  0.009402,   0.009402,    0.009402,    0.009402,
  0.009617,   0.009617,    0.009617,    0.009617,
  0.00981,    0.00981,     0.00981,     0.00981,
  0.01024,    0.01024,     0.01024,     0.01024,
  0.009756,   0.009756,    0.009756,    0.009756,
  0.008797,   0.008797,    0.008797,    0.008797,
  0.008608,   0.008608,    0.008608,    0.008608,
  0.008765,   0.008765,    0.008765,    0.008765,
  0.008829,   0.008829,    0.008829,    0.008829,
  0.008483,   0.008483,    0.008483,    0.008483,
  0.008074,   0.008074,    0.008074,    0.008074,
  0.0077,     0.0077,      0.0077,      0.0077,
  0.007388,   0.007388,    0.007388,    0.007388,
  0.00733,    0.00733,     0.00733,     0.00733,
  0.007395,   0.007395,    0.007395,    0.007395,
  0.00752,    0.00752,     0.00752,     0.00752,
  0.007671,   0.007671,    0.007671,    0.007671,
  0.007917,   0.007917,    0.007917,    0.007917,
  0.00798,    0.00798,     0.00798,     0.00798,
  0.007758,   0.007758,    0.007758,    0.007758,
  0.00779,    0.00779,     0.00779,     0.00779,
  0.007953,   0.007953,    0.007953,    0.007953,
  0.007965,   0.007965,    0.007965,    0.007965,
  0.008009,   0.008009,    0.008009,    0.008009,
  0.008055,   0.008055,    0.008055,    0.008055,
  0.00804,    0.00804,     0.00804,     0.00804,
  0.008008,   0.008008,    0.008008,    0.008008,
  0.007971,   0.007971,    0.007971,    0.007971,
  0.008019,   0.008019,    0.008019,    0.008019,
  0.008103,   0.008103,    0.008103,    0.008103,
  0.008157,   0.008157,    0.008157,    0.008157,
  0.008107,   0.008107,    0.008107,    0.008107,
  0.008006,   0.008006,    0.008006,    0.008006,
  0.00798,    0.00798,     0.00798,     0.00798,
  0.007894,   0.007894,    0.007894,    0.007894,
  0.007753,   0.007753,    0.007753,    0.007753,
  0.007624,   0.007624,    0.007624,    0.007624,
  0.007506,   0.007506,    0.007506,    0.007506,
  0.007436,   0.007436,    0.007436,    0.007436,
  0.007424,   0.007424,    0.007424,    0.007424,
  0.007446,   0.007446,    0.007446,    0.007446,
  0.007433,   0.007433,    0.007433,    0.007433,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.007575,   0.007575,    0.007575,    0.007575,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.008057,   0.008057,    0.008057,    0.008057,
  0.008563,   0.008563,    0.008563,    0.008563,
  0.008778,   0.008778,    0.008778,    0.008778,
  0.008868,   0.008868,    0.008868,    0.008868,
  0.008875,   0.008875,    0.008875,    0.008875,
  0.008656,   0.008656,    0.008656,    0.008656,
  0.008391,   0.008391,    0.008391,    0.008391,
  0.008139,   0.008139,    0.008139,    0.008139,
  0.00801,    0.00801,     0.00801,     0.00801,
  0.008076,   0.008076,    0.008076,    0.008076,
  0.007825,   0.007825,    0.007825,    0.007825,
  0.007015,   0.007015,    0.007015,    0.007015,
  0.0063,     0.0063,      0.0063,      0.0063,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.005798,   0.005798,    0.005798,    0.005798,
  0.00567,    0.00567,     0.00567,     0.00567,
  0.005855,   0.005855,    0.005855,    0.005855,
  0.006002,   0.006002,    0.006002,    0.006002,
  0.005932,   0.005932,    0.005932,    0.005932,
  0.005899,   0.005899,    0.005899,    0.005899,
  0.006026,   0.006026,    0.006026,    0.006026,
  0.00625,    0.00625,     0.00625,     0.00625,
  0.006555,   0.006555,    0.006555,    0.006555,
  0.006709,   0.006709,    0.006709,    0.006709,
  0.006742,   0.006742,    0.006742,    0.006742,
  0.006917,   0.006917,    0.006917,    0.006917,
  0.007105,   0.007105,    0.007105,    0.007105,
  0.007198,   0.007198,    0.007198,    0.007198,
  0.007246,   0.007246,    0.007246,    0.007246,
  0.007274,   0.007274,    0.007274,    0.007274,
  0.007386,   0.007386,    0.007386,    0.007386,
  0.007527,   0.007527,    0.007527,    0.007527,
  0.007647,   0.007647,    0.007647,    0.007647,
  0.007751,   0.007751,    0.007751,    0.007751,
  0.008077,   0.008077,    0.008077,    0.008077,
  0.008465,   0.008465,    0.008465,    0.008465,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.00853,    0.00853,     0.00853,     0.00853,
  0.00853,    0.00853,     0.00853,     0.00853,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.00853,    0.00853,     0.00853,     0.00853,
  0.00853,    0.00853,     0.00853,     0.00853,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.008579,   0.008579,    0.008579,    0.008579,
  0.008579,   0.008579,    0.008579,    0.008579,
  0.008579,   0.008579,    0.008579,    0.008579,
  0.008604,   0.008604,    0.008604,    0.008604,
  0.008678,   0.008678,    0.008678,    0.008678,
  0.008804,   0.008804,    0.008804,    0.008804,
  0.008905,   0.008905,    0.008905,    0.008905,
  0.009008,   0.009008,    0.009008,    0.009008,
  0.00919,    0.00919,     0.00919,     0.00919,
  0.00929,    0.00929,     0.00929,     0.00929,
  0.009419,   0.009419,    0.009419,    0.009419,
  0.009451,   0.009451,    0.009451,    0.009451,
  0.009232,   0.009232,    0.009232,    0.009232,
  0.00911,    0.00911,     0.00911,     0.00911,
  0.009139,   0.009139,    0.009139,    0.009139,
  0.009013,   0.009013,    0.009013,    0.009013,
  0.008515,   0.008515,    0.008515,    0.008515,
  0.008086,   0.008086,    0.008086,    0.008086,
  0.008085,   0.008085,    0.008085,    0.008085,
  0.008019,   0.008019,    0.008019,    0.008019,
  0.007763,   0.007763,    0.007763,    0.007763,
  0.007601,   0.007601,    0.007601,    0.007601,
  0.007569,   0.007569,    0.007569,    0.007569,
  0.007606,   0.007606,    0.007606,    0.007606,
  0.007675,   0.007675,    0.007675,    0.007675,
  0.007807,   0.007807,    0.007807,    0.007807,
  0.007923,   0.007923,    0.007923,    0.007923,
  0.007963,   0.007963,    0.007963,    0.007963,
  0.007949,   0.007949,    0.007949,    0.007949,
  0.00801,    0.00801,     0.00801,     0.00801,
  0.008119,   0.008119,    0.008119,    0.008119,
  0.008208,   0.008208,    0.008208,    0.008208,
  0.008278,   0.008278,    0.008278,    0.008278,
  0.008296,   0.008296,    0.008296,    0.008296,
  0.008306,   0.008306,    0.008306,    0.008306,
  0.008297,   0.008297,    0.008297,    0.008297,
  0.008328,   0.008328,    0.008328,    0.008328,
  0.00836,    0.00836,     0.00836,     0.00836,
  0.00836,    0.00836,     0.00836,     0.00836,
  0.008432,   0.008432,    0.008432,    0.008432,
  0.008506,   0.008506,    0.008506,    0.008506,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.008629,   0.008629,    0.008629,    0.008629,
  0.008703,   0.008703,    0.008703,    0.008703,
  0.008753,   0.008753,    0.008753,    0.008753,
  0.008804,   0.008804,    0.008804,    0.008804,
  0.008854,   0.008854,    0.008854,    0.008854,
  0.008905,   0.008905,    0.008905,    0.008905,
  0.008956,   0.008956,    0.008956,    0.008956,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.009008,   0.009008,    0.009008,    0.009008,
  0.009138,   0.009138,    0.009138,    0.009138,
  0.009281,   0.009281,    0.009281,    0.009281,
  0.009302,   0.009302,    0.009302,    0.009302,
  0.009267,   0.009267,    0.009267,    0.009267,
  0.009003,   0.009003,    0.009003,    0.009003,
  0.008625,   0.008625,    0.008625,    0.008625,
  0.008394,   0.008394,    0.008394,    0.008394,
  0.00817,    0.00817,     0.00817,     0.00817,
  0.007921,   0.007921,    0.007921,    0.007921,
  0.007582,   0.007582,    0.007582,    0.007582,
  0.007306,   0.007306,    0.007306,    0.007306,
  0.007306,   0.007306,    0.007306,    0.007306,
  0.007397,   0.007397,    0.007397,    0.007397,
  0.007424,   0.007424,    0.007424,    0.007424,
  0.007424,   0.007424,    0.007424,    0.007424,
  0.007364,   0.007364,    0.007364,    0.007364,
  0.007331,   0.007331,    0.007331,    0.007331,
  0.007427,   0.007427,    0.007427,    0.007427,
  0.00756,    0.00756,     0.00756,     0.00756,
  0.007759,   0.007759,    0.007759,    0.007759,
  0.007963,   0.007963,    0.007963,    0.007963,
  0.008043,   0.008043,    0.008043,    0.008043,
  0.008236,   0.008236,    0.008236,    0.008236,
  0.008519,   0.008519,    0.008519,    0.008519,
  0.008653,   0.008653,    0.008653,    0.008653,
  0.008658,   0.008658,    0.008658,    0.008658,
  0.008622,   0.008622,    0.008622,    0.008622,
  0.008617,   0.008617,    0.008617,    0.008617,
  0.008653,   0.008653,    0.008653,    0.008653,
  0.008694,   0.008694,    0.008694,    0.008694,
  0.008703,   0.008703,    0.008703,    0.008703,
  0.008708,   0.008708,    0.008708,    0.008708,
  0.008708,   0.008708,    0.008708,    0.008708,
  0.00866,    0.00866,     0.00866,     0.00866,
  0.008617,   0.008617,    0.008617,    0.008617,
  0.008654,   0.008654,    0.008654,    0.008654,
  0.008764,   0.008764,    0.008764,    0.008764,
  0.008801,   0.008801,    0.008801,    0.008801,
  0.008744,   0.008744,    0.008744,    0.008744,
  0.008685,   0.008685,    0.008685,    0.008685,
  0.008628,   0.008628,    0.008628,    0.008628,
  0.00859,    0.00859,     0.00859,     0.00859,
  0.008453,   0.008453,    0.008453,    0.008453,
  0.008261,   0.008261,    0.008261,    0.008261,
  0.008156,   0.008156,    0.008156,    0.008156,
  0.008117,   0.008117,    0.008117,    0.008117,
  0.008128,   0.008128,    0.008128,    0.008128,
  0.008188,   0.008188,    0.008188,    0.008188,
  0.008237,   0.008237,    0.008237,    0.008237,
  0.008252,   0.008252,    0.008252,    0.008252,
  0.008193,   0.008193,    0.008193,    0.008193,
  0.007984,   0.007984,    0.007984,    0.007984,
  0.007661,   0.007661,    0.007661,    0.007661,
  0.007258,   0.007258,    0.007258,    0.007258,
  0.007032,   0.007032,    0.007032,    0.007032,
  0.006985,   0.006985,    0.006985,    0.006985,
  0.006654,   0.006654,    0.006654,    0.006654,
  0.006173,   0.006173,    0.006173,    0.006173,
  0.005912,   0.005912,    0.005912,    0.005912,
  0.005688,   0.005688,    0.005688,    0.005688,
  0.005693,   0.005693,    0.005693,    0.005693,
  0.005729,   0.005729,    0.005729,    0.005729,
  0.005668,   0.005668,    0.005668,    0.005668,
  0.005894,   0.005894,    0.005894,    0.005894,
  0.006124,   0.006124,    0.006124,    0.006124,
  0.00634,    0.00634,     0.00634,     0.00634,
  0.006131,   0.006131,    0.006131,    0.006131,
  0.005764,   0.005764,    0.005764,    0.005764,
  0.005726,   0.005726,    0.005726,    0.005726,
  0.005486,   0.005486,    0.005486,    0.005486,
  0.005382,   0.005382,    0.005382,    0.005382,
  0.005715,   0.005715,    0.005715,    0.005715,
  0.006097,   0.006097,    0.006097,    0.006097,
  0.006265,   0.006265,    0.006265,    0.006265,
  0.006218,   0.006218,    0.006218,    0.006218,
  0.005895,   0.005895,    0.005895,    0.005895,
  0.005603,   0.005603,    0.005603,    0.005603,
  0.005626,   0.005626,    0.005626,    0.005626,
  0.005783,   0.005783,    0.005783,    0.005783,
  0.006012,   0.006012,    0.006012,    0.006012,
  0.006111,   0.006111,    0.006111,    0.006111,
  0.005726,   0.005726,    0.005726,    0.005726,
  0.005225,   0.005225,    0.005225,    0.005225,
  0.005059,   0.005059,    0.005059,    0.005059,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005164,   0.005164,    0.005164,    0.005164,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005567,   0.005567,    0.005567,    0.005567,
  0.005745,   0.005745,    0.005745,    0.005745,
  0.005855,   0.005855,    0.005855,    0.005855,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005884,   0.005884,    0.005884,    0.005884,
  0.005926,   0.005926,    0.005926,    0.005926,
  0.005957,   0.005957,    0.005957,    0.005957,
  0.005999,   0.005999,    0.005999,    0.005999,
  0.006031,   0.006031,    0.006031,    0.006031,
  0.006095,   0.006095,    0.006095,    0.006095,
  0.00613,    0.00613,     0.00613,     0.00613,
  0.006087,   0.006087,    0.006087,    0.006087,
  0.006004,   0.006004,    0.006004,    0.006004,
  0.005887,   0.005887,    0.005887,    0.005887,
  0.005682,   0.005682,    0.005682,    0.005682,
  0.005552,   0.005552,    0.005552,    0.005552,
  0.005478,   0.005478,    0.005478,    0.005478,
  0.005483,   0.005483,    0.005483,    0.005483,
  0.005464,   0.005464,    0.005464,    0.005464,
  0.005418,   0.005418,    0.005418,    0.005418,
  0.005409,   0.005409,    0.005409,    0.005409,
  0.005364,   0.005364,    0.005364,    0.005364,
  0.005439,   0.005439,    0.005439,    0.005439,
  0.005376,   0.005376,    0.005376,    0.005376,
  0.005302,   0.005302,    0.005302,    0.005302,
  0.005237,   0.005237,    0.005237,    0.005237,
  0.005159,   0.005159,    0.005159,    0.005159,
  0.005317,   0.005317,    0.005317,    0.005317,
  0.005629,   0.005629,    0.005629,    0.005629,
  0.005714,   0.005714,    0.005714,    0.005714,
  0.005624,   0.005624,    0.005624,    0.005624,
  0.005716,   0.005716,    0.005716,    0.005716,
  0.005879,   0.005879,    0.005879,    0.005879,
  0.005976,   0.005976,    0.005976,    0.005976,
  0.006009,   0.006009,    0.006009,    0.006009,
  0.0061,     0.0061,      0.0061,      0.0061,
  0.006194,   0.006194,    0.006194,    0.006194,
  0.006197,   0.006197,    0.006197,    0.006197,
  0.006156,   0.006156,    0.006156,    0.006156,
  0.006145,   0.006145,    0.006145,    0.006145,
  0.006161,   0.006161,    0.006161,    0.006161,
  0.00617,    0.00617,     0.00617,     0.00617,
  0.006169,   0.006169,    0.006169,    0.006169,
  0.006093,   0.006093,    0.006093,    0.006093,
  0.006064,   0.006064,    0.006064,    0.006064,
  0.00607,    0.00607,     0.00607,     0.00607,
  0.006026,   0.006026,    0.006026,    0.006026,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006076,   0.006076,    0.006076,    0.006076,
  0.006076,   0.006076,    0.006076,    0.006076,
  0.006102,   0.006102,    0.006102,    0.006102,
  0.006102,   0.006102,    0.006102,    0.006102,
  0.006044,   0.006044,    0.006044,    0.006044,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.006045,   0.006045,    0.006045,    0.006045,
  0.00607,    0.00607,     0.00607,     0.00607,
  0.006132,   0.006132,    0.006132,    0.006132,
  0.006275,   0.006275,    0.006275,    0.006275,
  0.006509,   0.006509,    0.006509,    0.006509,
  0.006645,   0.006645,    0.006645,    0.006645,
  0.006652,   0.006652,    0.006652,    0.006652,
  0.006402,   0.006402,    0.006402,    0.006402,
  0.006107,   0.006107,    0.006107,    0.006107,
  0.005963,   0.005963,    0.005963,    0.005963,
  0.005834,   0.005834,    0.005834,    0.005834,
  0.005767,   0.005767,    0.005767,    0.005767,
  0.005741,   0.005741,    0.005741,    0.005741,
  0.005729,   0.005729,    0.005729,    0.005729,
  0.005691,   0.005691,    0.005691,    0.005691,
  0.005652,   0.005652,    0.005652,    0.005652,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005553,   0.005553,    0.005553,    0.005553,
  0.005489,   0.005489,    0.005489,    0.005489,
  0.005553,   0.005553,    0.005553,    0.005553,
  0.005742,   0.005742,    0.005742,    0.005742,
  0.005964,   0.005964,    0.005964,    0.005964,
  0.006188,   0.006188,    0.006188,    0.006188,
  0.006473,   0.006473,    0.006473,    0.006473,
  0.006663,   0.006663,    0.006663,    0.006663,
  0.006831,   0.006831,    0.006831,    0.006831,
  0.006989,   0.006989,    0.006989,    0.006989,
  0.007134,   0.007134,    0.007134,    0.007134,
  0.007214,   0.007214,    0.007214,    0.007214,
  0.007212,   0.007212,    0.007212,    0.007212,
  0.007236,   0.007236,    0.007236,    0.007236,
  0.00721,    0.00721,     0.00721,     0.00721,
  0.007149,   0.007149,    0.007149,    0.007149,
  0.007138,   0.007138,    0.007138,    0.007138,
  0.007175,   0.007175,    0.007175,    0.007175,
  0.007242,   0.007242,    0.007242,    0.007242,
  0.007284,   0.007284,    0.007284,    0.007284,
  0.007368,   0.007368,    0.007368,    0.007368,
  0.007479,   0.007479,    0.007479,    0.007479,
  0.007547,   0.007547,    0.007547,    0.007547,
  0.007606,   0.007606,    0.007606,    0.007606,
  0.007654,   0.007654,    0.007654,    0.007654,
  0.007691,   0.007691,    0.007691,    0.007691,
  0.007773,   0.007773,    0.007773,    0.007773,
  0.008099,   0.008099,    0.008099,    0.008099,
  0.008484,   0.008484,    0.008484,    0.008484,
  0.008667,   0.008667,    0.008667,    0.008667,
  0.008796,   0.008796,    0.008796,    0.008796,
  0.008895,   0.008895,    0.008895,    0.008895,
  0.008975,   0.008975,    0.008975,    0.008975,
  0.009059,   0.009059,    0.009059,    0.009059,
  0.009131,   0.009131,    0.009131,    0.009131,
  0.009156,   0.009156,    0.009156,    0.009156,
  0.009001,   0.009001,    0.009001,    0.009001,
  0.008733,   0.008733,    0.008733,    0.008733,
  0.008472,   0.008472,    0.008472,    0.008472,
  0.008178,   0.008178,    0.008178,    0.008178,
  0.007845,   0.007845,    0.007845,    0.007845,
  0.007423,   0.007423,    0.007423,    0.007423,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007002,   0.007002,    0.007002,    0.007002,
  0.007004,   0.007004,    0.007004,    0.007004,
  0.007098,   0.007098,    0.007098,    0.007098,
  0.00716,    0.00716,     0.00716,     0.00716,
  0.00716,    0.00716,     0.00716,     0.00716,
  0.00719,    0.00719,     0.00719,     0.00719,
  0.007222,   0.007222,    0.007222,    0.007222,
  0.007224,   0.007224,    0.007224,    0.007224,
  0.007162,   0.007162,    0.007162,    0.007162,
  0.007131,   0.007131,    0.007131,    0.007131,
  0.007288,   0.007288,    0.007288,    0.007288,
  0.007445,   0.007445,    0.007445,    0.007445,
  0.007571,   0.007571,    0.007571,    0.007571,
  0.00773,    0.00773,     0.00773,     0.00773,
  0.007734,   0.007734,    0.007734,    0.007734,
  0.007676,   0.007676,    0.007676,    0.007676,
  0.008073,   0.008073,    0.008073,    0.008073,
  0.008484,   0.008484,    0.008484,    0.008484,
  0.008457,   0.008457,    0.008457,    0.008457,
  0.008258,   0.008258,    0.008258,    0.008258,
  0.008054,   0.008054,    0.008054,    0.008054,
  0.008045,   0.008045,    0.008045,    0.008045,
  0.008099,   0.008099,    0.008099,    0.008099,
  0.008067,   0.008067,    0.008067,    0.008067,
  0.008004,   0.008004,    0.008004,    0.008004,
  0.007928,   0.007928,    0.007928,    0.007928,
  0.007844,   0.007844,    0.007844,    0.007844,
  0.00789,    0.00789,     0.00789,     0.00789,
  0.008028,   0.008028,    0.008028,    0.008028,
  0.008005,   0.008005,    0.008005,    0.008005,
  0.007813,   0.007813,    0.007813,    0.007813,
  0.00769,    0.00769,     0.00769,     0.00769,
  0.007557,   0.007557,    0.007557,    0.007557,
  0.007274,   0.007274,    0.007274,    0.007274,
  0.006903,   0.006903,    0.006903,    0.006903,
  0.006632,   0.006632,    0.006632,    0.006632,
  0.006489,   0.006489,    0.006489,    0.006489,
  0.006405,   0.006405,    0.006405,    0.006405,
  0.006496,   0.006496,    0.006496,    0.006496,
  0.006695,   0.006695,    0.006695,    0.006695,
  0.006757,   0.006757,    0.006757,    0.006757,
  0.006651,   0.006651,    0.006651,    0.006651,
  0.006631,   0.006631,    0.006631,    0.006631,
  0.006641,   0.006641,    0.006641,    0.006641,
  0.006406,   0.006406,    0.006406,    0.006406,
  0.005937,   0.005937,    0.005937,    0.005937,
  0.005425,   0.005425,    0.005425,    0.005425,
  0.004938,   0.004938,    0.004938,    0.004938,
  0.004691,   0.004691,    0.004691,    0.004691,
  0.004701,   0.004701,    0.004701,    0.004701,
  0.004633,   0.004633,    0.004633,    0.004633,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004419,   0.004419,    0.004419,    0.004419,
  0.004172,   0.004172,    0.004172,    0.004172,
  0.004114,   0.004114,    0.004114,    0.004114,
  0.004204,   0.004204,    0.004204,    0.004204,
  0.004791,   0.004791,    0.004791,    0.004791,
  0.005649,   0.005649,    0.005649,    0.005649,
  0.006004,   0.006004,    0.006004,    0.006004,
  0.005823,   0.005823,    0.005823,    0.005823,
  0.005626,   0.005626,    0.005626,    0.005626,
  0.005605,   0.005605,    0.005605,    0.005605,
  0.005647,   0.005647,    0.005647,    0.005647,
  0.005603,   0.005603,    0.005603,    0.005603,
  0.005649,   0.005649,    0.005649,    0.005649,
  0.005699,   0.005699,    0.005699,    0.005699,
  0.005699,   0.005699,    0.005699,    0.005699,
  0.005787,   0.005787,    0.005787,    0.005787,
  0.005807,   0.005807,    0.005807,    0.005807,
  0.005803,   0.005803,    0.005803,    0.005803,
  0.006086,   0.006086,    0.006086,    0.006086,
  0.006389,   0.006389,    0.006389,    0.006389,
  0.006415,   0.006415,    0.006415,    0.006415,
  0.00634,    0.00634,     0.00634,     0.00634,
  0.006266,   0.006266,    0.006266,    0.006266,
  0.006191,   0.006191,    0.006191,    0.006191,
  0.006134,   0.006134,    0.006134,    0.006134,
  0.006134,   0.006134,    0.006134,    0.006134,
  0.006096,   0.006096,    0.006096,    0.006096,
  0.006014,   0.006014,    0.006014,    0.006014,
  0.006014,   0.006014,    0.006014,    0.006014,
  0.006022,   0.006022,    0.006022,    0.006022,
  0.005982,   0.005982,    0.005982,    0.005982,
  0.005895,   0.005895,    0.005895,    0.005895,
  0.005806,   0.005806,    0.005806,    0.005806,
  0.005819,   0.005819,    0.005819,    0.005819,
  0.005899,   0.005899,    0.005899,    0.005899,
  0.005994,   0.005994,    0.005994,    0.005994,
  0.006122,   0.006122,    0.006122,    0.006122,
  0.006246,   0.006246,    0.006246,    0.006246,
  0.006313,   0.006313,    0.006313,    0.006313,
  0.006306,   0.006306,    0.006306,    0.006306,
  0.006119,   0.006119,    0.006119,    0.006119,
  0.006108,   0.006108,    0.006108,    0.006108,
  0.005976,   0.005976,    0.005976,    0.005976,
  0.005467,   0.005467,    0.005467,    0.005467,
  0.005035,   0.005035,    0.005035,    0.005035,
  0.004893,   0.004893,    0.004893,    0.004893,
  0.004903,   0.004903,    0.004903,    0.004903,
  0.005021,   0.005021,    0.005021,    0.005021,
  0.00534,    0.00534,     0.00534,     0.00534,
  0.005502,   0.005502,    0.005502,    0.005502,
  0.005537,   0.005537,    0.005537,    0.005537,
  0.005456,   0.005456,    0.005456,    0.005456,
  0.00534,    0.00534,     0.00534,     0.00534,
  0.005354,   0.005354,    0.005354,    0.005354,
  0.005506,   0.005506,    0.005506,    0.005506,
  0.005756,   0.005756,    0.005756,    0.005756,
  0.005851,   0.005851,    0.005851,    0.005851,
  0.00588,    0.00588,     0.00588,     0.00588,
  0.006031,   0.006031,    0.006031,    0.006031,
  0.006163,   0.006163,    0.006163,    0.006163,
  0.006207,   0.006207,    0.006207,    0.006207,
  0.006183,   0.006183,    0.006183,    0.006183,
  0.006155,   0.006155,    0.006155,    0.006155,
  0.006117,   0.006117,    0.006117,    0.006117,
  0.006083,   0.006083,    0.006083,    0.006083,
  0.006104,   0.006104,    0.006104,    0.006104,
  0.006147,   0.006147,    0.006147,    0.006147,
  0.006172,   0.006172,    0.006172,    0.006172,
  0.006176,   0.006176,    0.006176,    0.006176,
  0.006179,   0.006179,    0.006179,    0.006179,
  0.006191,   0.006191,    0.006191,    0.006191,
  0.006262,   0.006262,    0.006262,    0.006262,
  0.006294,   0.006294,    0.006294,    0.006294,
  0.006266,   0.006266,    0.006266,    0.006266,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.006071,   0.006071,    0.006071,    0.006071,
  0.006115,   0.006115,    0.006115,    0.006115,
  0.006158,   0.006158,    0.006158,    0.006158,
  0.006183,   0.006183,    0.006183,    0.006183,
  0.006258,   0.006258,    0.006258,    0.006258,
  0.006413,   0.006413,    0.006413,    0.006413,
  0.006498,   0.006498,    0.006498,    0.006498,
  0.006523,   0.006523,    0.006523,    0.006523,
  0.006558,   0.006558,    0.006558,    0.006558,
  0.006563,   0.006563,    0.006563,    0.006563,
  0.006602,   0.006602,    0.006602,    0.006602,
  0.006654,   0.006654,    0.006654,    0.006654,
  0.006741,   0.006741,    0.006741,    0.006741,
  0.006686,   0.006686,    0.006686,    0.006686,
  0.006521,   0.006521,    0.006521,    0.006521,
  0.006435,   0.006435,    0.006435,    0.006435,
  0.006307,   0.006307,    0.006307,    0.006307,
  0.006179,   0.006179,    0.006179,    0.006179,
  0.006136,   0.006136,    0.006136,    0.006136,
  0.006065,   0.006065,    0.006065,    0.006065,
  0.005961,   0.005961,    0.005961,    0.005961,
  0.005826,   0.005826,    0.005826,    0.005826,
  0.00566,    0.00566,     0.00566,     0.00566,
  0.005566,   0.005566,    0.005566,    0.005566,
  0.00563,    0.00563,     0.00563,     0.00563,
  0.005626,   0.005626,    0.005626,    0.005626,
  0.005469,   0.005469,    0.005469,    0.005469,
  0.005539,   0.005539,    0.005539,    0.005539,
  0.005802,   0.005802,    0.005802,    0.005802,
  0.005979,   0.005979,    0.005979,    0.005979,
  0.006056,   0.006056,    0.006056,    0.006056,
  0.006169,   0.006169,    0.006169,    0.006169,
  0.006261,   0.006261,    0.006261,    0.006261,
  0.006305,   0.006305,    0.006305,    0.006305,
  0.006384,   0.006384,    0.006384,    0.006384,
  0.006436,   0.006436,    0.006436,    0.006436,
  0.006445,   0.006445,    0.006445,    0.006445,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.006458,   0.006458,    0.006458,    0.006458,
  0.006453,   0.006453,    0.006453,    0.006453,
  0.006408,   0.006408,    0.006408,    0.006408,
  0.00639,    0.00639,     0.00639,     0.00639,
  0.006387,   0.006387,    0.006387,    0.006387,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006282,   0.006282,    0.006282,    0.006282,
  0.006264,   0.006264,    0.006264,    0.006264,
  0.006279,   0.006279,    0.006279,    0.006279,
  0.006283,   0.006283,    0.006283,    0.006283,
  0.006315,   0.006315,    0.006315,    0.006315,
  0.006359,   0.006359,    0.006359,    0.006359,
  0.006349,   0.006349,    0.006349,    0.006349,
  0.006332,   0.006332,    0.006332,    0.006332,
  0.006302,   0.006302,    0.006302,    0.006302,
  0.006221,   0.006221,    0.006221,    0.006221,
  0.006195,   0.006195,    0.006195,    0.006195,
  0.006287,   0.006287,    0.006287,    0.006287,
  0.006395,   0.006395,    0.006395,    0.006395,
  0.006573,   0.006573,    0.006573,    0.006573,
  0.00689,    0.00689,     0.00689,     0.00689,
  0.007157,   0.007157,    0.007157,    0.007157,
  0.007311,   0.007311,    0.007311,    0.007311,
  0.006971,   0.006971,    0.006971,    0.006971,
  0.006434,   0.006434,    0.006434,    0.006434,
  0.006005,   0.006005,    0.006005,    0.006005,
  0.005521,   0.005521,    0.005521,    0.005521,
  0.00521,    0.00521,     0.00521,     0.00521,
  0.005002,   0.005002,    0.005002,    0.005002,
  0.004865,   0.004865,    0.004865,    0.004865,
  0.004791,   0.004791,    0.004791,    0.004791,
  0.004536,   0.004536,    0.004536,    0.004536,
  0.004212,   0.004212,    0.004212,    0.004212,
  0.004077,   0.004077,    0.004077,    0.004077,
  0.003949,   0.003949,    0.003949,    0.003949,
  0.004048,   0.004048,    0.004048,    0.004048,
  0.00437,    0.00437,     0.00437,     0.00437,
  0.004705,   0.004705,    0.004705,    0.004705,
  0.005096,   0.005096,    0.005096,    0.005096,
  0.0055,     0.0055,      0.0055,      0.0055,
  0.005807,   0.005807,    0.005807,    0.005807,
  0.006011,   0.006011,    0.006011,    0.006011,
  0.006194,   0.006194,    0.006194,    0.006194,
  0.006349,   0.006349,    0.006349,    0.006349,
  0.00638,    0.00638,     0.00638,     0.00638,
  0.006345,   0.006345,    0.006345,    0.006345,
  0.006368,   0.006368,    0.006368,    0.006368,
  0.006387,   0.006387,    0.006387,    0.006387,
  0.006392,   0.006392,    0.006392,    0.006392,
  0.006372,   0.006372,    0.006372,    0.006372,
  0.006373,   0.006373,    0.006373,    0.006373,
  0.0064,     0.0064,      0.0064,      0.0064,
  0.006515,   0.006515,    0.006515,    0.006515,
  0.006696,   0.006696,    0.006696,    0.006696,
  0.006827,   0.006827,    0.006827,    0.006827,
  0.006882,   0.006882,    0.006882,    0.006882,
  0.006902,   0.006902,    0.006902,    0.006902,
  0.006941,   0.006941,    0.006941,    0.006941,
  0.006964,   0.006964,    0.006964,    0.006964,
  0.006981,   0.006981,    0.006981,    0.006981,
  0.006991,   0.006991,    0.006991,    0.006991,
  0.006962,   0.006962,    0.006962,    0.006962,
  0.006948,   0.006948,    0.006948,    0.006948,
  0.006957,   0.006957,    0.006957,    0.006957,
  0.006925,   0.006925,    0.006925,    0.006925,
  0.006903,   0.006903,    0.006903,    0.006903,
  0.006963,   0.006963,    0.006963,    0.006963,
  0.007142,   0.007142,    0.007142,    0.007142,
  0.007364,   0.007364,    0.007364,    0.007364,
  0.007593,   0.007593,    0.007593,    0.007593,
  0.007823,   0.007823,    0.007823,    0.007823,
  0.007992,   0.007992,    0.007992,    0.007992,
  0.008151,   0.008151,    0.008151,    0.008151,
  0.008204,   0.008204,    0.008204,    0.008204,
  0.008172,   0.008172,    0.008172,    0.008172,
  0.008268,   0.008268,    0.008268,    0.008268,
  0.008457,   0.008457,    0.008457,    0.008457,
  0.008551,   0.008551,    0.008551,    0.008551,
  0.008518,   0.008518,    0.008518,    0.008518,
  0.008611,   0.008611,    0.008611,    0.008611,
  0.008673,   0.008673,    0.008673,    0.008673,
  0.008736,   0.008736,    0.008736,    0.008736,
  0.008994,   0.008994,    0.008994,    0.008994,
  0.009186,   0.009186,    0.009186,    0.009186,
  0.009316,   0.009316,    0.009316,    0.009316,
  0.009454,   0.009454,    0.009454,    0.009454,
  0.009552,   0.009552,    0.009552,    0.009552,
  0.009586,   0.009586,    0.009586,    0.009586,
  0.009625,   0.009625,    0.009625,    0.009625,
  0.009666,   0.009666,    0.009666,    0.009666,
  0.009646,   0.009646,    0.009646,    0.009646,
  0.009592,   0.009592,    0.009592,    0.009592,
  0.009568,   0.009568,    0.009568,    0.009568,
  0.009515,   0.009515,    0.009515,    0.009515,
  0.009376,   0.009376,    0.009376,    0.009376,
  0.009185,   0.009185,    0.009185,    0.009185,
  0.009007,   0.009007,    0.009007,    0.009007,
  0.008839,   0.008839,    0.008839,    0.008839,
  0.00864,    0.00864,     0.00864,     0.00864,
  0.008391,   0.008391,    0.008391,    0.008391,
  0.008171,   0.008171,    0.008171,    0.008171,
  0.008059,   0.008059,    0.008059,    0.008059,
  0.007981,   0.007981,    0.007981,    0.007981,
  0.007942,   0.007942,    0.007942,    0.007942,
  0.007927,   0.007927,    0.007927,    0.007927,
  0.007867,   0.007867,    0.007867,    0.007867,
  0.007776,   0.007776,    0.007776,    0.007776,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007641,   0.007641,    0.007641,    0.007641,
  0.007641,   0.007641,    0.007641,    0.007641,
  0.007641,   0.007641,    0.007641,    0.007641,
  0.007641,   0.007641,    0.007641,    0.007641,
  0.007709,   0.007709,    0.007709,    0.007709,
  0.007821,   0.007821,    0.007821,    0.007821,
  0.00803,    0.00803,     0.00803,     0.00803,
  0.008337,   0.008337,    0.008337,    0.008337,
  0.00868,    0.00868,     0.00868,     0.00868,
  0.009061,   0.009061,    0.009061,    0.009061,
  0.009161,   0.009161,    0.009161,    0.009161,
  0.008957,   0.008957,    0.008957,    0.008957,
  0.008821,   0.008821,    0.008821,    0.008821,
  0.008646,   0.008646,    0.008646,    0.008646,
  0.008576,   0.008576,    0.008576,    0.008576,
  0.008674,   0.008674,    0.008674,    0.008674,
  0.008563,   0.008563,    0.008563,    0.008563,
  0.008458,   0.008458,    0.008458,    0.008458,
  0.008474,   0.008474,    0.008474,    0.008474,
  0.008518,   0.008518,    0.008518,    0.008518,
  0.008521,   0.008521,    0.008521,    0.008521,
  0.008489,   0.008489,    0.008489,    0.008489,
  0.008641,   0.008641,    0.008641,    0.008641,
  0.008906,   0.008906,    0.008906,    0.008906,
  0.008954,   0.008954,    0.008954,    0.008954,
  0.008844,   0.008844,    0.008844,    0.008844,
  0.0088,     0.0088,      0.0088,      0.0088,
  0.008767,   0.008767,    0.008767,    0.008767,
  0.008784,   0.008784,    0.008784,    0.008784,
  0.008733,   0.008733,    0.008733,    0.008733,
  0.008544,   0.008544,    0.008544,    0.008544,
  0.008298,   0.008298,    0.008298,    0.008298,
  0.008043,   0.008043,    0.008043,    0.008043,
  0.007962,   0.007962,    0.007962,    0.007962,
  0.007928,   0.007928,    0.007928,    0.007928,
  0.007776,   0.007776,    0.007776,    0.007776,
  0.007642,   0.007642,    0.007642,    0.007642,
  0.007548,   0.007548,    0.007548,    0.007548,
  0.00747,    0.00747,     0.00747,     0.00747,
  0.007446,   0.007446,    0.007446,    0.007446,
  0.007382,   0.007382,    0.007382,    0.007382,
  0.007359,   0.007359,    0.007359,    0.007359,
  0.007398,   0.007398,    0.007398,    0.007398,
  0.007343,   0.007343,    0.007343,    0.007343,
  0.007303,   0.007303,    0.007303,    0.007303,
  0.007342,   0.007342,    0.007342,    0.007342,
  0.007335,   0.007335,    0.007335,    0.007335,
  0.00732,    0.00732,     0.00732,     0.00732,
  0.007291,   0.007291,    0.007291,    0.007291,
  0.007187,   0.007187,    0.007187,    0.007187,
  0.007106,   0.007106,    0.007106,    0.007106,
  0.007071,   0.007071,    0.007071,    0.007071,
  0.00703,    0.00703,     0.00703,     0.00703,
  0.007047,   0.007047,    0.007047,    0.007047,
  0.006994,   0.006994,    0.006994,    0.006994,
  0.006848,   0.006848,    0.006848,    0.006848,
  0.006665,   0.006665,    0.006665,    0.006665,
  0.006299,   0.006299,    0.006299,    0.006299,
  0.005914,   0.005914,    0.005914,    0.005914,
  0.005785,   0.005785,    0.005785,    0.005785,
  0.005846,   0.005846,    0.005846,    0.005846,
  0.00595,    0.00595,     0.00595,     0.00595,
  0.005951,   0.005951,    0.005951,    0.005951,
  0.005855,   0.005855,    0.005855,    0.005855,
  0.005758,   0.005758,    0.005758,    0.005758,
  0.005753,   0.005753,    0.005753,    0.005753,
  0.005913,   0.005913,    0.005913,    0.005913,
  0.00609,    0.00609,     0.00609,     0.00609,
  0.006085,   0.006085,    0.006085,    0.006085,
  0.005779,   0.005779,    0.005779,    0.005779,
  0.005428,   0.005428,    0.005428,    0.005428,
  0.00528,    0.00528,     0.00528,     0.00528,
  0.005177,   0.005177,    0.005177,    0.005177,
  0.004833,   0.004833,    0.004833,    0.004833,
  0.004438,   0.004438,    0.004438,    0.004438,
  0.004414,   0.004414,    0.004414,    0.004414,
  0.004604,   0.004604,    0.004604,    0.004604,
  0.004794,   0.004794,    0.004794,    0.004794,
  0.004977,   0.004977,    0.004977,    0.004977,
  0.005174,   0.005174,    0.005174,    0.005174,
  0.005359,   0.005359,    0.005359,    0.005359,
  0.005476,   0.005476,    0.005476,    0.005476,
  0.005604,   0.005604,    0.005604,    0.005604,
  0.005693,   0.005693,    0.005693,    0.005693,
  0.005711,   0.005711,    0.005711,    0.005711,
  0.005746,   0.005746,    0.005746,    0.005746,
  0.005763,   0.005763,    0.005763,    0.005763,
  0.005754,   0.005754,    0.005754,    0.005754,
  0.00573,    0.00573,     0.00573,     0.00573,
  0.005669,   0.005669,    0.005669,    0.005669,
  0.00565,    0.00565,     0.00565,     0.00565,
  0.005654,   0.005654,    0.005654,    0.005654,
  0.005623,   0.005623,    0.005623,    0.005623,
  0.00558,    0.00558,     0.00558,     0.00558,
  0.005542,   0.005542,    0.005542,    0.005542,
  0.005508,   0.005508,    0.005508,    0.005508,
  0.005388,   0.005388,    0.005388,    0.005388,
  0.005203,   0.005203,    0.005203,    0.005203,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005336,   0.005336,    0.005336,    0.005336,
  0.005772,   0.005772,    0.005772,    0.005772,
  0.006038,   0.006038,    0.006038,    0.006038,
  0.005983,   0.005983,    0.005983,    0.005983,
  0.005511,   0.005511,    0.005511,    0.005511,
  0.004936,   0.004936,    0.004936,    0.004936,
  0.004523,   0.004523,    0.004523,    0.004523,
  0.004338,   0.004338,    0.004338,    0.004338,
  0.004337,   0.004337,    0.004337,    0.004337,
  0.004269,   0.004269,    0.004269,    0.004269,
  0.004326,   0.004326,    0.004326,    0.004326,
  0.004501,   0.004501,    0.004501,    0.004501,
  0.004426,   0.004426,    0.004426,    0.004426,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.00425,    0.00425,     0.00425,     0.00425,
  0.004245,   0.004245,    0.004245,    0.004245,
  0.004267,   0.004267,    0.004267,    0.004267,
  0.004284,   0.004284,    0.004284,    0.004284,
  0.004199,   0.004199,    0.004199,    0.004199,
  0.004208,   0.004208,    0.004208,    0.004208,
  0.004351,   0.004351,    0.004351,    0.004351,
  0.004695,   0.004695,    0.004695,    0.004695,
  0.005107,   0.005107,    0.005107,    0.005107,
  0.005317,   0.005317,    0.005317,    0.005317,
  0.005368,   0.005368,    0.005368,    0.005368,
  0.005392,   0.005392,    0.005392,    0.005392,
  0.005394,   0.005394,    0.005394,    0.005394,
  0.005395,   0.005395,    0.005395,    0.005395,
  0.005373,   0.005373,    0.005373,    0.005373,
  0.005272,   0.005272,    0.005272,    0.005272,
  0.005258,   0.005258,    0.005258,    0.005258,
  0.005356,   0.005356,    0.005356,    0.005356,
  0.005404,   0.005404,    0.005404,    0.005404,
  0.005434,   0.005434,    0.005434,    0.005434,
  0.005515,   0.005515,    0.005515,    0.005515,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005601,   0.005601,    0.005601,    0.005601,
  0.005604,   0.005604,    0.005604,    0.005604,
  0.005596,   0.005596,    0.005596,    0.005596,
  0.005552,   0.005552,    0.005552,    0.005552,
  0.005545,   0.005545,    0.005545,    0.005545,
  0.005542,   0.005542,    0.005542,    0.005542,
  0.005525,   0.005525,    0.005525,    0.005525,
  0.005539,   0.005539,    0.005539,    0.005539,
  0.005536,   0.005536,    0.005536,    0.005536,
  0.005485,   0.005485,    0.005485,    0.005485,
  0.005468,   0.005468,    0.005468,    0.005468,
  0.005543,   0.005543,    0.005543,    0.005543,
  0.005675,   0.005675,    0.005675,    0.005675,
  0.005747,   0.005747,    0.005747,    0.005747,
  0.00571,    0.00571,     0.00571,     0.00571,
  0.005678,   0.005678,    0.005678,    0.005678,
  0.00568,    0.00568,     0.00568,     0.00568,
  0.00559,    0.00559,     0.00559,     0.00559,
  0.005364,   0.005364,    0.005364,    0.005364,
  0.005144,   0.005144,    0.005144,    0.005144,
  0.005018,   0.005018,    0.005018,    0.005018,
  0.005034,   0.005034,    0.005034,    0.005034,
  0.005058,   0.005058,    0.005058,    0.005058,
  0.005033,   0.005033,    0.005033,    0.005033,
  0.005067,   0.005067,    0.005067,    0.005067,
  0.005022,   0.005022,    0.005022,    0.005022,
  0.004978,   0.004978,    0.004978,    0.004978,
  0.005057,   0.005057,    0.005057,    0.005057,
  0.005084,   0.005084,    0.005084,    0.005084,
  0.005049,   0.005049,    0.005049,    0.005049,
  0.005018,   0.005018,    0.005018,    0.005018,
  0.005065,   0.005065,    0.005065,    0.005065,
  0.005121,   0.005121,    0.005121,    0.005121,
  0.005175,   0.005175,    0.005175,    0.005175,
  0.005392,   0.005392,    0.005392,    0.005392,
  0.005583,   0.005583,    0.005583,    0.005583,
  0.005607,   0.005607,    0.005607,    0.005607,
  0.005582,   0.005582,    0.005582,    0.005582,
  0.005572,   0.005572,    0.005572,    0.005572,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005523,   0.005523,    0.005523,    0.005523,
  0.005432,   0.005432,    0.005432,    0.005432,
  0.005392,   0.005392,    0.005392,    0.005392,
  0.005384,   0.005384,    0.005384,    0.005384,
  0.005392,   0.005392,    0.005392,    0.005392,
  0.005377,   0.005377,    0.005377,    0.005377,
  0.005357,   0.005357,    0.005357,    0.005357,
  0.00537,    0.00537,     0.00537,     0.00537,
  0.005402,   0.005402,    0.005402,    0.005402,
  0.005415,   0.005415,    0.005415,    0.005415,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005422,   0.005422,    0.005422,    0.005422,
  0.005425,   0.005425,    0.005425,    0.005425,
  0.005397,   0.005397,    0.005397,    0.005397,
  0.005371,   0.005371,    0.005371,    0.005371,
  0.00536,    0.00536,     0.00536,     0.00536,
  0.005367,   0.005367,    0.005367,    0.005367,
  0.005379,   0.005379,    0.005379,    0.005379,
  0.005438,   0.005438,    0.005438,    0.005438,
  0.005483,   0.005483,    0.005483,    0.005483,
  0.005457,   0.005457,    0.005457,    0.005457,
  0.005448,   0.005448,    0.005448,    0.005448,
  0.005437,   0.005437,    0.005437,    0.005437,
  0.005339,   0.005339,    0.005339,    0.005339,
  0.005155,   0.005155,    0.005155,    0.005155,
  0.004976,   0.004976,    0.004976,    0.004976,
  0.00492,    0.00492,     0.00492,     0.00492,
  0.005011,   0.005011,    0.005011,    0.005011,
  0.005142,   0.005142,    0.005142,    0.005142,
  0.005213,   0.005213,    0.005213,    0.005213,
  0.005163,   0.005163,    0.005163,    0.005163,
  0.004963,   0.004963,    0.004963,    0.004963,
  0.004861,   0.004861,    0.004861,    0.004861,
  0.004923,   0.004923,    0.004923,    0.004923,
  0.004986,   0.004986,    0.004986,    0.004986,
  0.005049,   0.005049,    0.005049,    0.005049,
  0.005111,   0.005111,    0.005111,    0.005111,
  0.005206,   0.005206,    0.005206,    0.005206,
  0.005241,   0.005241,    0.005241,    0.005241,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005659,   0.005659,    0.005659,    0.005659,
  0.005974,   0.005974,    0.005974,    0.005974,
  0.006158,   0.006158,    0.006158,    0.006158,
  0.00625,    0.00625,     0.00625,     0.00625,
  0.006281,   0.006281,    0.006281,    0.006281,
  0.006241,   0.006241,    0.006241,    0.006241,
  0.006233,   0.006233,    0.006233,    0.006233,
  0.006323,   0.006323,    0.006323,    0.006323,
  0.006431,   0.006431,    0.006431,    0.006431,
  0.006515,   0.006515,    0.006515,    0.006515,
  0.006536,   0.006536,    0.006536,    0.006536,
  0.006518,   0.006518,    0.006518,    0.006518,
  0.0065,     0.0065,      0.0065,      0.0065,
  0.006509,   0.006509,    0.006509,    0.006509,
  0.006548,   0.006548,    0.006548,    0.006548,
  0.006557,   0.006557,    0.006557,    0.006557,
  0.006548,   0.006548,    0.006548,    0.006548,
  0.006529,   0.006529,    0.006529,    0.006529,
  0.00646,    0.00646,     0.00646,     0.00646,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006278,   0.006278,    0.006278,    0.006278,
  0.006208,   0.006208,    0.006208,    0.006208,
  0.006171,   0.006171,    0.006171,    0.006171,
  0.006152,   0.006152,    0.006152,    0.006152,
  0.006128,   0.006128,    0.006128,    0.006128,
  0.006104,   0.006104,    0.006104,    0.006104,
  0.006184,   0.006184,    0.006184,    0.006184,
  0.006328,   0.006328,    0.006328,    0.006328,
  0.006558,   0.006558,    0.006558,    0.006558,
  0.006863,   0.006863,    0.006863,    0.006863,
  0.006986,   0.006986,    0.006986,    0.006986,
  0.006982,   0.006982,    0.006982,    0.006982,
  0.006885,   0.006885,    0.006885,    0.006885,
  0.006675,   0.006675,    0.006675,    0.006675,
  0.006395,   0.006395,    0.006395,    0.006395,
  0.006108,   0.006108,    0.006108,    0.006108,
  0.006029,   0.006029,    0.006029,    0.006029,
  0.005917,   0.005917,    0.005917,    0.005917,
  0.005798,   0.005798,    0.005798,    0.005798,
  0.005813,   0.005813,    0.005813,    0.005813,
  0.005835,   0.005835,    0.005835,    0.005835,
  0.005926,   0.005926,    0.005926,    0.005926,
  0.006155,   0.006155,    0.006155,    0.006155,
  0.006529,   0.006529,    0.006529,    0.006529,
  0.006916,   0.006916,    0.006916,    0.006916,
  0.007083,   0.007083,    0.007083,    0.007083,
  0.00708,    0.00708,     0.00708,     0.00708,
  0.007131,   0.007131,    0.007131,    0.007131,
  0.007184,   0.007184,    0.007184,    0.007184,
  0.007181,   0.007181,    0.007181,    0.007181,
  0.007191,   0.007191,    0.007191,    0.007191,
  0.007219,   0.007219,    0.007219,    0.007219,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007243,   0.007243,    0.007243,    0.007243,
  0.007257,   0.007257,    0.007257,    0.007257,
  0.00732,    0.00732,     0.00732,     0.00732,
  0.007407,   0.007407,    0.007407,    0.007407,
  0.007446,   0.007446,    0.007446,    0.007446,
  0.0075,     0.0075,      0.0075,      0.0075,
  0.007518,   0.007518,    0.007518,    0.007518,
  0.007426,   0.007426,    0.007426,    0.007426,
  0.007339,   0.007339,    0.007339,    0.007339,
  0.007282,   0.007282,    0.007282,    0.007282,
  0.007186,   0.007186,    0.007186,    0.007186,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007292,   0.007292,    0.007292,    0.007292,
  0.007378,   0.007378,    0.007378,    0.007378,
  0.007465,   0.007465,    0.007465,    0.007465,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007531,   0.007531,    0.007531,    0.007531,
  0.007597,   0.007597,    0.007597,    0.007597,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007822,   0.007822,    0.007822,    0.007822,
  0.00799,    0.00799,     0.00799,     0.00799,
  0.008141,   0.008141,    0.008141,    0.008141,
  0.008213,   0.008213,    0.008213,    0.008213,
  0.008156,   0.008156,    0.008156,    0.008156,
  0.008109,   0.008109,    0.008109,    0.008109,
  0.008161,   0.008161,    0.008161,    0.008161,
  0.008159,   0.008159,    0.008159,    0.008159,
  0.008069,   0.008069,    0.008069,    0.008069,
  0.007935,   0.007935,    0.007935,    0.007935,
  0.007766,   0.007766,    0.007766,    0.007766,
  0.007618,   0.007618,    0.007618,    0.007618,
  0.007485,   0.007485,    0.007485,    0.007485,
  0.007391,   0.007391,    0.007391,    0.007391,
  0.007331,   0.007331,    0.007331,    0.007331,
  0.007369,   0.007369,    0.007369,    0.007369,
  0.007499,   0.007499,    0.007499,    0.007499,
  0.007506,   0.007506,    0.007506,    0.007506,
  0.00753,    0.00753,     0.00753,     0.00753,
  0.007677,   0.007677,    0.007677,    0.007677,
  0.007754,   0.007754,    0.007754,    0.007754,
  0.007804,   0.007804,    0.007804,    0.007804,
  0.00783,    0.00783,     0.00783,     0.00783,
  0.007762,   0.007762,    0.007762,    0.007762,
  0.007659,   0.007659,    0.007659,    0.007659,
  0.007626,   0.007626,    0.007626,    0.007626,
  0.007639,   0.007639,    0.007639,    0.007639,
  0.007575,   0.007575,    0.007575,    0.007575,
  0.007448,   0.007448,    0.007448,    0.007448,
  0.007297,   0.007297,    0.007297,    0.007297,
  0.007137,   0.007137,    0.007137,    0.007137,
  0.007018,   0.007018,    0.007018,    0.007018,
  0.006913,   0.006913,    0.006913,    0.006913,
  0.006841,   0.006841,    0.006841,    0.006841,
  0.006811,   0.006811,    0.006811,    0.006811,
  0.006811,   0.006811,    0.006811,    0.006811,
  0.00682,    0.00682,     0.00682,     0.00682,
  0.006798,   0.006798,    0.006798,    0.006798,
  0.006787,   0.006787,    0.006787,    0.006787,
  0.006798,   0.006798,    0.006798,    0.006798,
  0.006841,   0.006841,    0.006841,    0.006841,
  0.006861,   0.006861,    0.006861,    0.006861,
  0.00685,    0.00685,     0.00685,     0.00685,
  0.006809,   0.006809,    0.006809,    0.006809,
  0.006768,   0.006768,    0.006768,    0.006768,
  0.006707,   0.006707,    0.006707,    0.006707,
  0.006626,   0.006626,    0.006626,    0.006626,
  0.006738,   0.006738,    0.006738,    0.006738,
  0.006995,   0.006995,    0.006995,    0.006995,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007155,   0.007155,    0.007155,    0.007155,
  0.007114,   0.007114,    0.007114,    0.007114,
  0.006795,   0.006795,    0.006795,    0.006795,
  0.006266,   0.006266,    0.006266,    0.006266,
  0.005965,   0.005965,    0.005965,    0.005965,
  0.005774,   0.005774,    0.005774,    0.005774,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005571,   0.005571,    0.005571,    0.005571,
  0.005674,   0.005674,    0.005674,    0.005674,
  0.005802,   0.005802,    0.005802,    0.005802,
  0.005746,   0.005746,    0.005746,    0.005746,
  0.005475,   0.005475,    0.005475,    0.005475,
  0.005421,   0.005421,    0.005421,    0.005421,
  0.005456,   0.005456,    0.005456,    0.005456,
  0.005364,   0.005364,    0.005364,    0.005364,
  0.005327,   0.005327,    0.005327,    0.005327,
  0.005467,   0.005467,    0.005467,    0.005467,
  0.00592,    0.00592,     0.00592,     0.00592,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.006801,   0.006801,    0.006801,    0.006801,
  0.006959,   0.006959,    0.006959,    0.006959,
  0.006923,   0.006923,    0.006923,    0.006923,
  0.006782,   0.006782,    0.006782,    0.006782,
  0.006721,   0.006721,    0.006721,    0.006721,
  0.006807,   0.006807,    0.006807,    0.006807,
  0.006907,   0.006907,    0.006907,    0.006907,
  0.006872,   0.006872,    0.006872,    0.006872,
  0.006722,   0.006722,    0.006722,    0.006722,
  0.006593,   0.006593,    0.006593,    0.006593,
  0.006585,   0.006585,    0.006585,    0.006585,
  0.00665,    0.00665,     0.00665,     0.00665,
  0.006691,   0.006691,    0.006691,    0.006691,
  0.006697,   0.006697,    0.006697,    0.006697,
  0.006684,   0.006684,    0.006684,    0.006684,
  0.006687,   0.006687,    0.006687,    0.006687,
  0.006715,   0.006715,    0.006715,    0.006715,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006766,   0.006766,    0.006766,    0.006766,
  0.006725,   0.006725,    0.006725,    0.006725,
  0.006584,   0.006584,    0.006584,    0.006584,
  0.006549,   0.006549,    0.006549,    0.006549,
  0.006553,   0.006553,    0.006553,    0.006553,
  0.006507,   0.006507,    0.006507,    0.006507,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.006538,   0.006538,    0.006538,    0.006538,
  0.006703,   0.006703,    0.006703,    0.006703,
  0.006834,   0.006834,    0.006834,    0.006834,
  0.006828,   0.006828,    0.006828,    0.006828,
  0.006793,   0.006793,    0.006793,    0.006793,
  0.006835,   0.006835,    0.006835,    0.006835,
  0.007011,   0.007011,    0.007011,    0.007011,
  0.007089,   0.007089,    0.007089,    0.007089,
  0.007099,   0.007099,    0.007099,    0.007099,
  0.007203,   0.007203,    0.007203,    0.007203,
  0.007106,   0.007106,    0.007106,    0.007106,
  0.00691,    0.00691,     0.00691,     0.00691,
  0.007015,   0.007015,    0.007015,    0.007015,
  0.007152,   0.007152,    0.007152,    0.007152,
  0.007072,   0.007072,    0.007072,    0.007072,
  0.006804,   0.006804,    0.006804,    0.006804,
  0.006593,   0.006593,    0.006593,    0.006593,
  0.006564,   0.006564,    0.006564,    0.006564,
  0.006744,   0.006744,    0.006744,    0.006744,
  0.007164,   0.007164,    0.007164,    0.007164,
  0.007364,   0.007364,    0.007364,    0.007364,
  0.007446,   0.007446,    0.007446,    0.007446,
  0.007668,   0.007668,    0.007668,    0.007668,
  0.007877,   0.007877,    0.007877,    0.007877,
  0.008039,   0.008039,    0.008039,    0.008039,
  0.008168,   0.008168,    0.008168,    0.008168,
  0.008188,   0.008188,    0.008188,    0.008188,
  0.008094,   0.008094,    0.008094,    0.008094,
  0.007929,   0.007929,    0.007929,    0.007929,
  0.007753,   0.007753,    0.007753,    0.007753,
  0.007653,   0.007653,    0.007653,    0.007653,
  0.007587,   0.007587,    0.007587,    0.007587,
  0.007497,   0.007497,    0.007497,    0.007497,
  0.007439,   0.007439,    0.007439,    0.007439,
  0.007392,   0.007392,    0.007392,    0.007392,
  0.007294,   0.007294,    0.007294,    0.007294,
  0.007239,   0.007239,    0.007239,    0.007239,
  0.007335,   0.007335,    0.007335,    0.007335,
  0.007465,   0.007465,    0.007465,    0.007465,
  0.007477,   0.007477,    0.007477,    0.007477,
  0.007414,   0.007414,    0.007414,    0.007414,
  0.00732,    0.00732,     0.00732,     0.00732,
  0.007247,   0.007247,    0.007247,    0.007247,
  0.007238,   0.007238,    0.007238,    0.007238,
  0.007238,   0.007238,    0.007238,    0.007238,
  0.007216,   0.007216,    0.007216,    0.007216,
  0.007216,   0.007216,    0.007216,    0.007216,
  0.007238,   0.007238,    0.007238,    0.007238,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007232,   0.007232,    0.007232,    0.007232,
  0.007227,   0.007227,    0.007227,    0.007227,
  0.0072,     0.0072,      0.0072,      0.0072,
  0.007169,   0.007169,    0.007169,    0.007169,
  0.007177,   0.007177,    0.007177,    0.007177,
  0.007232,   0.007232,    0.007232,    0.007232,
  0.007246,   0.007246,    0.007246,    0.007246,
  0.007237,   0.007237,    0.007237,    0.007237,
  0.007205,   0.007205,    0.007205,    0.007205,
  0.007157,   0.007157,    0.007157,    0.007157,
  0.007107,   0.007107,    0.007107,    0.007107,
  0.007068,   0.007068,    0.007068,    0.007068,
  0.007051,   0.007051,    0.007051,    0.007051,
  0.006997,   0.006997,    0.006997,    0.006997,
  0.006959,   0.006959,    0.006959,    0.006959,
  0.006949,   0.006949,    0.006949,    0.006949,
  0.00693,    0.00693,     0.00693,     0.00693,
  0.00693,    0.00693,     0.00693,     0.00693,
  0.007002,   0.007002,    0.007002,    0.007002,
  0.007148,   0.007148,    0.007148,    0.007148,
  0.007273,   0.007273,    0.007273,    0.007273,
  0.007307,   0.007307,    0.007307,    0.007307,
  0.007351,   0.007351,    0.007351,    0.007351,
  0.007472,   0.007472,    0.007472,    0.007472,
  0.007453,   0.007453,    0.007453,    0.007453,
  0.007258,   0.007258,    0.007258,    0.007258,
  0.007082,   0.007082,    0.007082,    0.007082,
  0.006955,   0.006955,    0.006955,    0.006955,
  0.006841,   0.006841,    0.006841,    0.006841,
  0.006741,   0.006741,    0.006741,    0.006741,
  0.006624,   0.006624,    0.006624,    0.006624,
  0.006442,   0.006442,    0.006442,    0.006442,
  0.00618,    0.00618,     0.00618,     0.00618,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.005818,   0.005818,    0.005818,    0.005818,
  0.005629,   0.005629,    0.005629,    0.005629,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005249,   0.005249,    0.005249,    0.005249,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005249,   0.005249,    0.005249,    0.005249,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005395,   0.005395,    0.005395,    0.005395,
  0.005595,   0.005595,    0.005595,    0.005595,
  0.005855,   0.005855,    0.005855,    0.005855,
  0.006105,   0.006105,    0.006105,    0.006105,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.0065,     0.0065,      0.0065,      0.0065,
  0.006756,   0.006756,    0.006756,    0.006756,
  0.007234,   0.007234,    0.007234,    0.007234,
  0.007944,   0.007944,    0.007944,    0.007944,
  0.007842,   0.007842,    0.007842,    0.007842,
  0.007282,   0.007282,    0.007282,    0.007282,
  0.006984,   0.006984,    0.006984,    0.006984,
  0.006807,   0.006807,    0.006807,    0.006807,
  0.006889,   0.006889,    0.006889,    0.006889,
  0.006886,   0.006886,    0.006886,    0.006886,
  0.006917,   0.006917,    0.006917,    0.006917,
  0.007237,   0.007237,    0.007237,    0.007237,
  0.007603,   0.007603,    0.007603,    0.007603,
  0.007701,   0.007701,    0.007701,    0.007701,
  0.007725,   0.007725,    0.007725,    0.007725,
  0.007754,   0.007754,    0.007754,    0.007754,
  0.007715,   0.007715,    0.007715,    0.007715,
  0.007729,   0.007729,    0.007729,    0.007729,
  0.007779,   0.007779,    0.007779,    0.007779,
  0.00776,    0.00776,     0.00776,     0.00776,
  0.00763,    0.00763,     0.00763,     0.00763,
  0.007463,   0.007463,    0.007463,    0.007463,
  0.007304,   0.007304,    0.007304,    0.007304,
  0.006961,   0.006961,    0.006961,    0.006961,
  0.006755,   0.006755,    0.006755,    0.006755,
  0.006657,   0.006657,    0.006657,    0.006657,
  0.006133,   0.006133,    0.006133,    0.006133,
  0.005836,   0.005836,    0.005836,    0.005836,
  0.005717,   0.005717,    0.005717,    0.005717,
  0.005363,   0.005363,    0.005363,    0.005363,
  0.005154,   0.005154,    0.005154,    0.005154,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.004967,   0.004967,    0.004967,    0.004967,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005186,   0.005186,    0.005186,    0.005186,
  0.005497,   0.005497,    0.005497,    0.005497,
  0.005909,   0.005909,    0.005909,    0.005909,
  0.00637,    0.00637,     0.00637,     0.00637,
  0.006879,   0.006879,    0.006879,    0.006879,
  0.007294,   0.007294,    0.007294,    0.007294,
  0.007598,   0.007598,    0.007598,    0.007598,
  0.007891,   0.007891,    0.007891,    0.007891,
  0.008315,   0.008315,    0.008315,    0.008315,
  0.008275,   0.008275,    0.008275,    0.008275,
  0.00794,    0.00794,     0.00794,     0.00794,
  0.007892,   0.007892,    0.007892,    0.007892,
  0.007842,   0.007842,    0.007842,    0.007842,
  0.007804,   0.007804,    0.007804,    0.007804,
  0.007815,   0.007815,    0.007815,    0.007815,
  0.007771,   0.007771,    0.007771,    0.007771,
  0.007774,   0.007774,    0.007774,    0.007774,
  0.007865,   0.007865,    0.007865,    0.007865,
  0.007931,   0.007931,    0.007931,    0.007931,
  0.008,      0.008,       0.008,       0.008,
  0.008068,   0.008068,    0.008068,    0.008068,
  0.008056,   0.008056,    0.008056,    0.008056,
  0.007951,   0.007951,    0.007951,    0.007951,
  0.007944,   0.007944,    0.007944,    0.007944,
  0.00812,    0.00812,     0.00812,     0.00812,
  0.008287,   0.008287,    0.008287,    0.008287,
  0.008361,   0.008361,    0.008361,    0.008361,
  0.008424,   0.008424,    0.008424,    0.008424,
  0.008435,   0.008435,    0.008435,    0.008435,
  0.008446,   0.008446,    0.008446,    0.008446,
  0.008464,   0.008464,    0.008464,    0.008464,
  0.008389,   0.008389,    0.008389,    0.008389,
  0.008352,   0.008352,    0.008352,    0.008352,
  0.008377,   0.008377,    0.008377,    0.008377,
  0.008352,   0.008352,    0.008352,    0.008352,
  0.00831,    0.00831,     0.00831,     0.00831,
  0.008292,   0.008292,    0.008292,    0.008292,
  0.008324,   0.008324,    0.008324,    0.008324,
  0.008362,   0.008362,    0.008362,    0.008362,
  0.008425,   0.008425,    0.008425,    0.008425,
  0.008506,   0.008506,    0.008506,    0.008506,
  0.00853,    0.00853,     0.00853,     0.00853,
  0.00853,    0.00853,     0.00853,     0.00853,
  0.008555,   0.008555,    0.008555,    0.008555,
  0.008604,   0.008604,    0.008604,    0.008604,
  0.008653,   0.008653,    0.008653,    0.008653,
  0.008678,   0.008678,    0.008678,    0.008678,
  0.008678,   0.008678,    0.008678,    0.008678,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008855,   0.008855,    0.008855,    0.008855,
  0.009008,   0.009008,    0.009008,    0.009008,
  0.009163,   0.009163,    0.009163,    0.009163,
  0.009295,   0.009295,    0.009295,    0.009295,
  0.009401,   0.009401,    0.009401,    0.009401,
  0.009492,   0.009492,    0.009492,    0.009492,
  0.009377,   0.009377,    0.009377,    0.009377,
  0.008991,   0.008991,    0.008991,    0.008991,
  0.008749,   0.008749,    0.008749,    0.008749,
  0.008616,   0.008616,    0.008616,    0.008616,
  0.00836,    0.00836,     0.00836,     0.00836,
  0.008199,   0.008199,    0.008199,    0.008199,
  0.008104,   0.008104,    0.008104,    0.008104,
  0.00801,    0.00801,     0.00801,     0.00801,
  0.008011,   0.008011,    0.008011,    0.008011,
  0.008074,   0.008074,    0.008074,    0.008074,
  0.008073,   0.008073,    0.008073,    0.008073,
  0.008104,   0.008104,    0.008104,    0.008104,
  0.00839,    0.00839,     0.00839,     0.00839,
  0.008619,   0.008619,    0.008619,    0.008619,
  0.008661,   0.008661,    0.008661,    0.008661,
  0.008707,   0.008707,    0.008707,    0.008707,
  0.008779,   0.008779,    0.008779,    0.008779,
  0.009225,   0.009225,    0.009225,    0.009225,
  0.009712,   0.009712,    0.009712,    0.009712,
  0.009827,   0.009827,    0.009827,    0.009827,
  0.009619,   0.009619,    0.009619,    0.009619,
  0.009217,   0.009217,    0.009217,    0.009217,
  0.008956,   0.008956,    0.008956,    0.008956,
  0.008829,   0.008829,    0.008829,    0.008829,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008653,   0.008653,    0.008653,    0.008653,
  0.008629,   0.008629,    0.008629,    0.008629,
  0.008653,   0.008653,    0.008653,    0.008653,
  0.008678,   0.008678,    0.008678,    0.008678,
  0.008678,   0.008678,    0.008678,    0.008678,
  0.008703,   0.008703,    0.008703,    0.008703,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008728,   0.008728,    0.008728,    0.008728,
  0.008753,   0.008753,    0.008753,    0.008753,
  0.008778,   0.008778,    0.008778,    0.008778,
  0.008804,   0.008804,    0.008804,    0.008804,
  0.008854,   0.008854,    0.008854,    0.008854,
  0.00888,    0.00888,     0.00888,     0.00888,
  0.008931,   0.008931,    0.008931,    0.008931,
  0.009086,   0.009086,    0.009086,    0.009086,
  0.009349,   0.009349,    0.009349,    0.009349,
  0.009645,   0.009645,    0.009645,    0.009645,
  0.009893,   0.009893,    0.009893,    0.009893,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.0102,     0.0102,      0.0102,      0.0102,
  0.01032,    0.01032,     0.01032,     0.01032,
  0.01047,    0.01047,     0.01047,     0.01047,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01047,    0.01047,     0.01047,     0.01047,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01058,    0.01058,     0.01058,     0.01058,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01038,    0.01038,     0.01038,     0.01038,
  0.01044,    0.01044,     0.01044,     0.01044,
  0.01043,    0.01043,     0.01043,     0.01043,
  0.01027,    0.01027,     0.01027,     0.01027,
  0.01022,    0.01022,     0.01022,     0.01022,
  0.01025,    0.01025,     0.01025,     0.01025,
  0.0103,     0.0103,      0.0103,      0.0103,
  0.01033,    0.01033,     0.01033,     0.01033,
  0.01033,    0.01033,     0.01033,     0.01033,
  0.01033,    0.01033,     0.01033,     0.01033,
  0.0102,     0.0102,      0.0102,      0.0102,
  0.009987,   0.009987,    0.009987,    0.009987,
  0.009802,   0.009802,    0.009802,    0.009802,
  0.009681,   0.009681,    0.009681,    0.009681,
  0.009659,   0.009659,    0.009659,    0.009659,
  0.009455,   0.009455,    0.009455,    0.009455,
  0.009123,   0.009123,    0.009123,    0.009123,
  0.008834,   0.008834,    0.008834,    0.008834,
  0.008357,   0.008357,    0.008357,    0.008357,
  0.008091,   0.008091,    0.008091,    0.008091,
  0.007979,   0.007979,    0.007979,    0.007979,
  0.007773,   0.007773,    0.007773,    0.007773,
  0.007667,   0.007667,    0.007667,    0.007667,
  0.007562,   0.007562,    0.007562,    0.007562,
  0.007395,   0.007395,    0.007395,    0.007395,
  0.007261,   0.007261,    0.007261,    0.007261,
  0.00721,    0.00721,     0.00721,     0.00721,
  0.007153,   0.007153,    0.007153,    0.007153,
  0.007041,   0.007041,    0.007041,    0.007041,
  0.006906,   0.006906,    0.006906,    0.006906,
  0.006794,   0.006794,    0.006794,    0.006794,
  0.006787,   0.006787,    0.006787,    0.006787,
  0.006899,   0.006899,    0.006899,    0.006899,
  0.006917,   0.006917,    0.006917,    0.006917,
  0.006815,   0.006815,    0.006815,    0.006815,
  0.006777,   0.006777,    0.006777,    0.006777,
  0.006713,   0.006713,    0.006713,    0.006713,
  0.006466,   0.006466,    0.006466,    0.006466,
  0.00634,    0.00634,     0.00634,     0.00634,
  0.006114,   0.006114,    0.006114,    0.006114,
  0.006073,   0.006073,    0.006073,    0.006073,
  0.006281,   0.006281,    0.006281,    0.006281,
  0.006267,   0.006267,    0.006267,    0.006267,
  0.006301,   0.006301,    0.006301,    0.006301,
  0.005733,   0.005733,    0.005733,    0.005733,
  0.005116,   0.005116,    0.005116,    0.005116,
  0.005131,   0.005131,    0.005131,    0.005131,
  0.004876,   0.004876,    0.004876,    0.004876,
  0.00454,    0.00454,     0.00454,     0.00454,
  0.00478,    0.00478,     0.00478,     0.00478,
  0.005385,   0.005385,    0.005385,    0.005385,
  0.005952,   0.005952,    0.005952,    0.005952,
  0.006313,   0.006313,    0.006313,    0.006313,
  0.006485,   0.006485,    0.006485,    0.006485,
  0.006454,   0.006454,    0.006454,    0.006454,
  0.006224,   0.006224,    0.006224,    0.006224,
  0.006052,   0.006052,    0.006052,    0.006052,
  0.006058,   0.006058,    0.006058,    0.006058,
  0.006164,   0.006164,    0.006164,    0.006164,
  0.006244,   0.006244,    0.006244,    0.006244,
  0.006242,   0.006242,    0.006242,    0.006242,
  0.00621,    0.00621,     0.00621,     0.00621,
  0.006094,   0.006094,    0.006094,    0.006094,
  0.0058,     0.0058,      0.0058,      0.0058,
  0.005548,   0.005548,    0.005548,    0.005548,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005622,   0.005622,    0.005622,    0.005622,
  0.005666,   0.005666,    0.005666,    0.005666,
  0.005658,   0.005658,    0.005658,    0.005658,
  0.005661,   0.005661,    0.005661,    0.005661,
  0.005616,   0.005616,    0.005616,    0.005616,
  0.005541,   0.005541,    0.005541,    0.005541,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.00547,    0.00547,     0.00547,     0.00547,
  0.005451,   0.005451,    0.005451,    0.005451,
  0.005433,   0.005433,    0.005433,    0.005433,
  0.005438,   0.005438,    0.005438,    0.005438,
  0.005426,   0.005426,    0.005426,    0.005426,
  0.005399,   0.005399,    0.005399,    0.005399,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005399,   0.005399,    0.005399,    0.005399,
  0.00543,    0.00543,     0.00543,     0.00543,
  0.005462,   0.005462,    0.005462,    0.005462,
  0.005549,   0.005549,    0.005549,    0.005549,
  0.005761,   0.005761,    0.005761,    0.005761,
  0.005959,   0.005959,    0.005959,    0.005959,
  0.006039,   0.006039,    0.006039,    0.006039,
  0.006073,   0.006073,    0.006073,    0.006073,
  0.006243,   0.006243,    0.006243,    0.006243,
  0.0065,     0.0065,      0.0065,      0.0065,
  0.006675,   0.006675,    0.006675,    0.006675,
  0.006763,   0.006763,    0.006763,    0.006763,
  0.006914,   0.006914,    0.006914,    0.006914,
  0.007015,   0.007015,    0.007015,    0.007015,
  0.006919,   0.006919,    0.006919,    0.006919,
  0.006785,   0.006785,    0.006785,    0.006785,
  0.006712,   0.006712,    0.006712,    0.006712,
  0.006628,   0.006628,    0.006628,    0.006628,
  0.006612,   0.006612,    0.006612,    0.006612,
  0.006818,   0.006818,    0.006818,    0.006818,
  0.007009,   0.007009,    0.007009,    0.007009,
  0.007021,   0.007021,    0.007021,    0.007021,
  0.00699,    0.00699,     0.00699,     0.00699,
  0.007011,   0.007011,    0.007011,    0.007011,
  0.006994,   0.006994,    0.006994,    0.006994,
  0.006899,   0.006899,    0.006899,    0.006899,
  0.006833,   0.006833,    0.006833,    0.006833,
  0.006887,   0.006887,    0.006887,    0.006887,
  0.007043,   0.007043,    0.007043,    0.007043,
  0.007156,   0.007156,    0.007156,    0.007156,
  0.007178,   0.007178,    0.007178,    0.007178,
  0.007195,   0.007195,    0.007195,    0.007195,
  0.007174,   0.007174,    0.007174,    0.007174,
  0.007146,   0.007146,    0.007146,    0.007146,
  0.007145,   0.007145,    0.007145,    0.007145,
  0.007153,   0.007153,    0.007153,    0.007153,
  0.007208,   0.007208,    0.007208,    0.007208,
  0.007279,   0.007279,    0.007279,    0.007279,
  0.007342,   0.007342,    0.007342,    0.007342,
  0.00746,    0.00746,     0.00746,     0.00746,
  0.007578,   0.007578,    0.007578,    0.007578,
  0.007595,   0.007595,    0.007595,    0.007595,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007383,   0.007383,    0.007383,    0.007383,
  0.007296,   0.007296,    0.007296,    0.007296,
  0.007233,   0.007233,    0.007233,    0.007233,
  0.007219,   0.007219,    0.007219,    0.007219,
  0.00726,    0.00726,     0.00726,     0.00726,
  0.007323,   0.007323,    0.007323,    0.007323,
  0.007369,   0.007369,    0.007369,    0.007369,
  0.007407,   0.007407,    0.007407,    0.007407,
  0.007519,   0.007519,    0.007519,    0.007519,
  0.007624,   0.007624,    0.007624,    0.007624,
  0.007709,   0.007709,    0.007709,    0.007709,
  0.007845,   0.007845,    0.007845,    0.007845,
  0.007972,   0.007972,    0.007972,    0.007972,
  0.008073,   0.008073,    0.008073,    0.008073,
  0.008024,   0.008024,    0.008024,    0.008024,
  0.007986,   0.007986,    0.007986,    0.007986,
  0.007822,   0.007822,    0.007822,    0.007822,
  0.007501,   0.007501,    0.007501,    0.007501,
  0.007464,   0.007464,    0.007464,    0.007464,
  0.00753,    0.00753,     0.00753,     0.00753,
  0.007504,   0.007504,    0.007504,    0.007504,
  0.007507,   0.007507,    0.007507,    0.007507,
  0.007573,   0.007573,    0.007573,    0.007573,
  0.007545,   0.007545,    0.007545,    0.007545,
  0.007618,   0.007618,    0.007618,    0.007618,
  0.007877,   0.007877,    0.007877,    0.007877,
  0.007943,   0.007943,    0.007943,    0.007943,
  0.007825,   0.007825,    0.007825,    0.007825,
  0.007675,   0.007675,    0.007675,    0.007675,
  0.007601,   0.007601,    0.007601,    0.007601,
  0.007591,   0.007591,    0.007591,    0.007591,
  0.007589,   0.007589,    0.007589,    0.007589,
  0.007554,   0.007554,    0.007554,    0.007554,
  0.007481,   0.007481,    0.007481,    0.007481,
  0.007464,   0.007464,    0.007464,    0.007464,
  0.007505,   0.007505,    0.007505,    0.007505,
  0.007541,   0.007541,    0.007541,    0.007541,
  0.007492,   0.007492,    0.007492,    0.007492,
  0.007444,   0.007444,    0.007444,    0.007444,
  0.007405,   0.007405,    0.007405,    0.007405,
  0.007381,   0.007381,    0.007381,    0.007381,
  0.00746,    0.00746,     0.00746,     0.00746,
  0.007579,   0.007579,    0.007579,    0.007579,
  0.007667,   0.007667,    0.007667,    0.007667,
  0.007747,   0.007747,    0.007747,    0.007747,
  0.007818,   0.007818,    0.007818,    0.007818,
  0.007881,   0.007881,    0.007881,    0.007881,
  0.007982,   0.007982,    0.007982,    0.007982,
  0.008122,   0.008122,    0.008122,    0.008122,
  0.008216,   0.008216,    0.008216,    0.008216,
  0.008216,   0.008216,    0.008216,    0.008216,
  0.008169,   0.008169,    0.008169,    0.008169,
  0.008145,   0.008145,    0.008145,    0.008145,
  0.008193,   0.008193,    0.008193,    0.008193,
  0.008216,   0.008216,    0.008216,    0.008216,
  0.008169,   0.008169,    0.008169,    0.008169,
  0.008145,   0.008145,    0.008145,    0.008145,
  0.008122,   0.008122,    0.008122,    0.008122,
  0.008098,   0.008098,    0.008098,    0.008098,
  0.008145,   0.008145,    0.008145,    0.008145,
  0.008193,   0.008193,    0.008193,    0.008193,
  0.008216,   0.008216,    0.008216,    0.008216,
  0.008312,   0.008312,    0.008312,    0.008312,
  0.008457,   0.008457,    0.008457,    0.008457,
  0.008642,   0.008642,    0.008642,    0.008642,
  0.008777,   0.008777,    0.008777,    0.008777,
  0.008768,   0.008768,    0.008768,    0.008768,
  0.008652,   0.008652,    0.008652,    0.008652,
  0.008538,   0.008538,    0.008538,    0.008538,
  0.00851,    0.00851,     0.00851,     0.00851,
  0.008451,   0.008451,    0.008451,    0.008451,
  0.008168,   0.008168,    0.008168,    0.008168,
  0.007955,   0.007955,    0.007955,    0.007955,
  0.007971,   0.007971,    0.007971,    0.007971,
  0.007965,   0.007965,    0.007965,    0.007965,
  0.007993,   0.007993,    0.007993,    0.007993,
  0.00805,    0.00805,     0.00805,     0.00805,
  0.008109,   0.008109,    0.008109,    0.008109,
  0.008157,   0.008157,    0.008157,    0.008157,
  0.008137,   0.008137,    0.008137,    0.008137,
  0.008061,   0.008061,    0.008061,    0.008061,
  0.007991,   0.007991,    0.007991,    0.007991,
  0.007979,   0.007979,    0.007979,    0.007979,
  0.007992,   0.007992,    0.007992,    0.007992,
  0.007974,   0.007974,    0.007974,    0.007974,
  0.007949,   0.007949,    0.007949,    0.007949,
  0.007981,   0.007981,    0.007981,    0.007981,
  0.008019,   0.008019,    0.008019,    0.008019,
  0.008026,   0.008026,    0.008026,    0.008026,
  0.008002,   0.008002,    0.008002,    0.008002,
  0.007977,   0.007977,    0.007977,    0.007977,
  0.007928,   0.007928,    0.007928,    0.007928,
  0.00788,    0.00788,     0.00788,     0.00788,
  0.0078,     0.0078,      0.0078,      0.0078,
  0.007649,   0.007649,    0.007649,    0.007649,
  0.007579,   0.007579,    0.007579,    0.007579,
  0.007485,   0.007485,    0.007485,    0.007485,
  0.007299,   0.007299,    0.007299,    0.007299,
  0.007113,   0.007113,    0.007113,    0.007113,
  0.006967,   0.006967,    0.006967,    0.006967,
  0.006896,   0.006896,    0.006896,    0.006896,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006783,   0.006783,    0.006783,    0.006783,
  0.006792,   0.006792,    0.006792,    0.006792,
  0.006936,   0.006936,    0.006936,    0.006936,
  0.007128,   0.007128,    0.007128,    0.007128,
  0.007393,   0.007393,    0.007393,    0.007393,
  0.007602,   0.007602,    0.007602,    0.007602,
  0.007621,   0.007621,    0.007621,    0.007621,
  0.00753,    0.00753,     0.00753,     0.00753,
  0.007374,   0.007374,    0.007374,    0.007374,
  0.007159,   0.007159,    0.007159,    0.007159,
  0.006979,   0.006979,    0.006979,    0.006979,
  0.007035,   0.007035,    0.007035,    0.007035,
  0.007254,   0.007254,    0.007254,    0.007254,
  0.007352,   0.007352,    0.007352,    0.007352,
  0.00727,    0.00727,     0.00727,     0.00727,
  0.007241,   0.007241,    0.007241,    0.007241,
  0.007366,   0.007366,    0.007366,    0.007366,
  0.007438,   0.007438,    0.007438,    0.007438,
  0.007544,   0.007544,    0.007544,    0.007544,
  0.007727,   0.007727,    0.007727,    0.007727,
  0.007929,   0.007929,    0.007929,    0.007929,
  0.00817,    0.00817,     0.00817,     0.00817,
  0.008357,   0.008357,    0.008357,    0.008357,
  0.008359,   0.008359,    0.008359,    0.008359,
  0.008296,   0.008296,    0.008296,    0.008296,
  0.008296,   0.008296,    0.008296,    0.008296,
  0.008361,   0.008361,    0.008361,    0.008361,
  0.008492,   0.008492,    0.008492,    0.008492,
  0.008628,   0.008628,    0.008628,    0.008628,
  0.008733,   0.008733,    0.008733,    0.008733,
  0.00884,    0.00884,     0.00884,     0.00884,
  0.008916,   0.008916,    0.008916,    0.008916,
  0.008982,   0.008982,    0.008982,    0.008982,
  0.009036,   0.009036,    0.009036,    0.009036,
  0.009024,   0.009024,    0.009024,    0.009024,
  0.009009,   0.009009,    0.009009,    0.009009,
  0.009032,   0.009032,    0.009032,    0.009032,
  0.009284,   0.009284,    0.009284,    0.009284,
  0.009812,   0.009812,    0.009812,    0.009812,
  0.01006,    0.01006,     0.01006,     0.01006,
  0.009949,   0.009949,    0.009949,    0.009949,
  0.009865,   0.009865,    0.009865,    0.009865,
  0.009809,   0.009809,    0.009809,    0.009809,
  0.009782,   0.009782,    0.009782,    0.009782,
  0.009809,   0.009809,    0.009809,    0.009809,
  0.009837,   0.009837,    0.009837,    0.009837,
  0.009837,   0.009837,    0.009837,    0.009837,
  0.009865,   0.009865,    0.009865,    0.009865,
  0.009921,   0.009921,    0.009921,    0.009921,
  0.009949,   0.009949,    0.009949,    0.009949,
  0.009946,   0.009946,    0.009946,    0.009946,
  0.009974,   0.009974,    0.009974,    0.009974,
  0.01003,    0.01003,     0.01003,     0.01003,
  0.01005,    0.01005,     0.01005,     0.01005,
  0.01007,    0.01007,     0.01007,     0.01007,
  0.01011,    0.01011,     0.01011,     0.01011,
  0.01004,    0.01004,     0.01004,     0.01004,
  0.009714,   0.009714,    0.009714,    0.009714,
  0.009307,   0.009307,    0.009307,    0.009307,
  0.008939,   0.008939,    0.008939,    0.008939,
  0.008572,   0.008572,    0.008572,    0.008572,
  0.00827,    0.00827,     0.00827,     0.00827,
  0.008075,   0.008075,    0.008075,    0.008075,
  0.007997,   0.007997,    0.007997,    0.007997,
  0.007615,   0.007615,    0.007615,    0.007615,
  0.007399,   0.007399,    0.007399,    0.007399,
  0.007745,   0.007745,    0.007745,    0.007745,
  0.008014,   0.008014,    0.008014,    0.008014,
  0.008002,   0.008002,    0.008002,    0.008002,
  0.007876,   0.007876,    0.007876,    0.007876,
  0.007827,   0.007827,    0.007827,    0.007827,
  0.007802,   0.007802,    0.007802,    0.007802,
  0.007827,   0.007827,    0.007827,    0.007827,
  0.007648,   0.007648,    0.007648,    0.007648,
  0.00734,    0.00734,     0.00734,     0.00734,
  0.007134,   0.007134,    0.007134,    0.007134,
  0.006959,   0.006959,    0.006959,    0.006959,
  0.006902,   0.006902,    0.006902,    0.006902,
  0.006972,   0.006972,    0.006972,    0.006972,
  0.00698,    0.00698,     0.00698,     0.00698,
  0.006917,   0.006917,    0.006917,    0.006917,
  0.006878,   0.006878,    0.006878,    0.006878,
  0.006862,   0.006862,    0.006862,    0.006862,
  0.006901,   0.006901,    0.006901,    0.006901,
  0.006925,   0.006925,    0.006925,    0.006925,
  0.006848,   0.006848,    0.006848,    0.006848,
  0.00673,    0.00673,     0.00673,     0.00673,
  0.006627,   0.006627,    0.006627,    0.006627,
  0.006573,   0.006573,    0.006573,    0.006573,
  0.006548,   0.006548,    0.006548,    0.006548,
  0.006531,   0.006531,    0.006531,    0.006531,
  0.006563,   0.006563,    0.006563,    0.006563,
  0.006626,   0.006626,    0.006626,    0.006626,
  0.006744,   0.006744,    0.006744,    0.006744,
  0.006848,   0.006848,    0.006848,    0.006848,
  0.006966,   0.006966,    0.006966,    0.006966,
  0.0071,     0.0071,      0.0071,      0.0071,
  0.007156,   0.007156,    0.007156,    0.007156,
  0.007232,   0.007232,    0.007232,    0.007232,
  0.007286,   0.007286,    0.007286,    0.007286,
  0.007454,   0.007454,    0.007454,    0.007454,
  0.007816,   0.007816,    0.007816,    0.007816,
  0.008122,   0.008122,    0.008122,    0.008122,
  0.008361,   0.008361,    0.008361,    0.008361,
  0.00863,    0.00863,     0.00863,     0.00863,
  0.008932,   0.008932,    0.008932,    0.008932,
  0.009127,   0.009127,    0.009127,    0.009127,
  0.009275,   0.009275,    0.009275,    0.009275,
  0.009468,   0.009468,    0.009468,    0.009468,
  0.009636,   0.009636,    0.009636,    0.009636,
  0.009767,   0.009767,    0.009767,    0.009767,
  0.009816,   0.009816,    0.009816,    0.009816,
  0.00987,    0.00987,     0.00987,     0.00987,
  0.009887,   0.009887,    0.009887,    0.009887,
  0.009818,   0.009818,    0.009818,    0.009818,
  0.009773,   0.009773,    0.009773,    0.009773,
  0.009739,   0.009739,    0.009739,    0.009739,
  0.009687,   0.009687,    0.009687,    0.009687,
  0.009542,   0.009542,    0.009542,    0.009542,
  0.009414,   0.009414,    0.009414,    0.009414,
  0.009401,   0.009401,    0.009401,    0.009401,
  0.009455,   0.009455,    0.009455,    0.009455,
  0.009563,   0.009563,    0.009563,    0.009563,
  0.009644,   0.009644,    0.009644,    0.009644,
  0.009727,   0.009727,    0.009727,    0.009727,
  0.009893,   0.009893,    0.009893,    0.009893,
  0.01009,    0.01009,     0.01009,     0.01009,
  0.01029,    0.01029,     0.01029,     0.01029,
  0.01043,    0.01043,     0.01043,     0.01043,
  0.01045,    0.01045,     0.01045,     0.01045,
  0.01041,    0.01041,     0.01041,     0.01041,
  0.01035,    0.01035,     0.01035,     0.01035,
  0.01029,    0.01029,     0.01029,     0.01029,
  0.01026,    0.01026,     0.01026,     0.01026,
  0.01029,    0.01029,     0.01029,     0.01029,
  0.01042,    0.01042,     0.01042,     0.01042,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.01055,    0.01055,     0.01055,     0.01055,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01058,    0.01058,     0.01058,     0.01058,
  0.01061,    0.01061,     0.01061,     0.01061,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01047,    0.01047,     0.01047,     0.01047,
  0.01047,    0.01047,     0.01047,     0.01047,
  0.01052,    0.01052,     0.01052,     0.01052,
  0.01064,    0.01064,     0.01064,     0.01064,
  0.0107,     0.0107,      0.0107,      0.0107,
  0.0106,     0.0106,      0.0106,      0.0106,
  0.009965,   0.009965,    0.009965,    0.009965,
  0.009209,   0.009209,    0.009209,    0.009209,
  0.008893,   0.008893,    0.008893,    0.008893,
  0.008736,   0.008736,    0.008736,    0.008736,
  0.008769,   0.008769,    0.008769,    0.008769,
  0.008801,   0.008801,    0.008801,    0.008801,
  0.008673,   0.008673,    0.008673,    0.008673,
  0.008972,   0.008972,    0.008972,    0.008972,
  0.009436,   0.009436,    0.009436,    0.009436,
  0.009232,   0.009232,    0.009232,    0.009232,
  0.008895,   0.008895,    0.008895,    0.008895,
  0.008862,   0.008862,    0.008862,    0.008862,
  0.008832,   0.008832,    0.008832,    0.008832,
  0.008865,   0.008865,    0.008865,    0.008865,
  0.008963,   0.008963,    0.008963,    0.008963,
  0.008998,   0.008998,    0.008998,    0.008998,
  0.008939,   0.008939,    0.008939,    0.008939,
  0.008881,   0.008881,    0.008881,    0.008881,
  0.008944,   0.008944,    0.008944,    0.008944,
  0.008977,   0.008977,    0.008977,    0.008977,
  0.009022,   0.009022,    0.009022,    0.009022,
  0.009011,   0.009011,    0.009011,    0.009011,
  0.008903,   0.008903,    0.008903,    0.008903,
  0.008857,   0.008857,    0.008857,    0.008857,
  0.008813,   0.008813,    0.008813,    0.008813,
  0.008798,   0.008798,    0.008798,    0.008798,
  0.008842,   0.008842,    0.008842,    0.008842,
  0.008964,   0.008964,    0.008964,    0.008964,
  0.009077,   0.009077,    0.009077,    0.009077,
  0.00916,    0.00916,     0.00916,     0.00916,
  0.009207,   0.009207,    0.009207,    0.009207,
  0.009314,   0.009314,    0.009314,    0.009314,
  0.009459,   0.009459,    0.009459,    0.009459,
  0.009518,   0.009518,    0.009518,    0.009518,
  0.009514,   0.009514,    0.009514,    0.009514,
  0.009459,   0.009459,    0.009459,    0.009459,
  0.009468,   0.009468,    0.009468,    0.009468,
  0.009504,   0.009504,    0.009504,    0.009504,
  0.009508,   0.009508,    0.009508,    0.009508,
  0.009428,   0.009428,    0.009428,    0.009428,
  0.009348,   0.009348,    0.009348,    0.009348,
  0.009237,   0.009237,    0.009237,    0.009237,
  0.009132,   0.009132,    0.009132,    0.009132,
  0.009189,   0.009189,    0.009189,    0.009189,
  0.009179,   0.009179,    0.009179,    0.009179,
  0.009021,   0.009021,    0.009021,    0.009021,
  0.008922,   0.008922,    0.008922,    0.008922,
  0.008512,   0.008512,    0.008512,    0.008512,
  0.007643,   0.007643,    0.007643,    0.007643,
  0.007053,   0.007053,    0.007053,    0.007053,
  0.00672,    0.00672,     0.00672,     0.00672,
  0.00633,    0.00633,     0.00633,     0.00633,
  0.006084,   0.006084,    0.006084,    0.006084,
  0.006021,   0.006021,    0.006021,    0.006021,
  0.006004,   0.006004,    0.006004,    0.006004,
  0.00603,    0.00603,     0.00603,     0.00603,
  0.00611,    0.00611,     0.00611,     0.00611,
  0.006104,   0.006104,    0.006104,    0.006104,
  0.005998,   0.005998,    0.005998,    0.005998,
  0.005925,   0.005925,    0.005925,    0.005925,
  0.005956,   0.005956,    0.005956,    0.005956,
  0.005967,   0.005967,    0.005967,    0.005967,
  0.005941,   0.005941,    0.005941,    0.005941,
  0.006002,   0.006002,    0.006002,    0.006002,
  0.005962,   0.005962,    0.005962,    0.005962,
  0.005831,   0.005831,    0.005831,    0.005831,
  0.006183,   0.006183,    0.006183,    0.006183,
  0.006661,   0.006661,    0.006661,    0.006661,
  0.006777,   0.006777,    0.006777,    0.006777,
  0.006832,   0.006832,    0.006832,    0.006832,
  0.006734,   0.006734,    0.006734,    0.006734,
  0.006532,   0.006532,    0.006532,    0.006532,
  0.006554,   0.006554,    0.006554,    0.006554,
  0.006741,   0.006741,    0.006741,    0.006741,
  0.006935,   0.006935,    0.006935,    0.006935,
  0.007113,   0.007113,    0.007113,    0.007113,
  0.007188,   0.007188,    0.007188,    0.007188,
  0.007221,   0.007221,    0.007221,    0.007221,
  0.007252,   0.007252,    0.007252,    0.007252,
  0.007241,   0.007241,    0.007241,    0.007241,
  0.00725,    0.00725,     0.00725,     0.00725,
  0.00725,    0.00725,     0.00725,     0.00725,
  0.007239,   0.007239,    0.007239,    0.007239,
  0.007271,   0.007271,    0.007271,    0.007271,
  0.007306,   0.007306,    0.007306,    0.007306,
  0.00731,    0.00731,     0.00731,     0.00731,
  0.007269,   0.007269,    0.007269,    0.007269,
  0.007206,   0.007206,    0.007206,    0.007206,
  0.007143,   0.007143,    0.007143,    0.007143,
  0.007112,   0.007112,    0.007112,    0.007112,
  0.007036,   0.007036,    0.007036,    0.007036,
  0.006929,   0.006929,    0.006929,    0.006929,
  0.00691,    0.00691,     0.00691,     0.00691,
  0.006913,   0.006913,    0.006913,    0.006913,
  0.006986,   0.006986,    0.006986,    0.006986,
  0.007096,   0.007096,    0.007096,    0.007096,
  0.007155,   0.007155,    0.007155,    0.007155,
  0.007229,   0.007229,    0.007229,    0.007229,
  0.007252,   0.007252,    0.007252,    0.007252,
  0.007266,   0.007266,    0.007266,    0.007266,
  0.007101,   0.007101,    0.007101,    0.007101,
  0.006659,   0.006659,    0.006659,    0.006659,
  0.006357,   0.006357,    0.006357,    0.006357,
  0.006255,   0.006255,    0.006255,    0.006255,
  0.006179,   0.006179,    0.006179,    0.006179,
  0.006133,   0.006133,    0.006133,    0.006133,
  0.006133,   0.006133,    0.006133,    0.006133,
  0.006218,   0.006218,    0.006218,    0.006218,
  0.006408,   0.006408,    0.006408,    0.006408,
  0.006566,   0.006566,    0.006566,    0.006566,
  0.006693,   0.006693,    0.006693,    0.006693,
  0.00681,    0.00681,     0.00681,     0.00681,
  0.006724,   0.006724,    0.006724,    0.006724,
  0.00657,    0.00657,     0.00657,     0.00657,
  0.006697,   0.006697,    0.006697,    0.006697,
  0.006867,   0.006867,    0.006867,    0.006867,
  0.006904,   0.006904,    0.006904,    0.006904,
  0.006924,   0.006924,    0.006924,    0.006924,
  0.006923,   0.006923,    0.006923,    0.006923,
  0.006955,   0.006955,    0.006955,    0.006955,
  0.006956,   0.006956,    0.006956,    0.006956,
  0.006926,   0.006926,    0.006926,    0.006926,
  0.006876,   0.006876,    0.006876,    0.006876,
  0.006795,   0.006795,    0.006795,    0.006795,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006715,   0.006715,    0.006715,    0.006715,
  0.006695,   0.006695,    0.006695,    0.006695,
  0.006675,   0.006675,    0.006675,    0.006675,
  0.006675,   0.006675,    0.006675,    0.006675,
  0.006655,   0.006655,    0.006655,    0.006655,
  0.006596,   0.006596,    0.006596,    0.006596,
  0.006461,   0.006461,    0.006461,    0.006461,
  0.006272,   0.006272,    0.006272,    0.006272,
  0.006051,   0.006051,    0.006051,    0.006051,
  0.005854,   0.005854,    0.005854,    0.005854,
  0.005766,   0.005766,    0.005766,    0.005766,
  0.00568,    0.00568,     0.00568,     0.00568,
  0.005561,   0.005561,    0.005561,    0.005561,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005753,   0.005753,    0.005753,    0.005753,
  0.006316,   0.006316,    0.006316,    0.006316,
  0.006879,   0.006879,    0.006879,    0.006879,
  0.007184,   0.007184,    0.007184,    0.007184,
  0.007089,   0.007089,    0.007089,    0.007089,
  0.006919,   0.006919,    0.006919,    0.006919,
  0.006579,   0.006579,    0.006579,    0.006579,
  0.006313,   0.006313,    0.006313,    0.006313,
  0.006536,   0.006536,    0.006536,    0.006536,
  0.006263,   0.006263,    0.006263,    0.006263,
  0.005293,   0.005293,    0.005293,    0.005293,
  0.004666,   0.004666,    0.004666,    0.004666,
  0.004715,   0.004715,    0.004715,    0.004715,
  0.005173,   0.005173,    0.005173,    0.005173,
  0.005825,   0.005825,    0.005825,    0.005825,
  0.006088,   0.006088,    0.006088,    0.006088,
  0.005888,   0.005888,    0.005888,    0.005888,
  0.005667,   0.005667,    0.005667,    0.005667,
  0.005518,   0.005518,    0.005518,    0.005518,
  0.005466,   0.005466,    0.005466,    0.005466,
  0.005772,   0.005772,    0.005772,    0.005772,
  0.006121,   0.006121,    0.006121,    0.006121,
  0.006158,   0.006158,    0.006158,    0.006158,
  0.006171,   0.006171,    0.006171,    0.006171,
  0.006176,   0.006176,    0.006176,    0.006176,
  0.006189,   0.006189,    0.006189,    0.006189,
  0.006208,   0.006208,    0.006208,    0.006208,
  0.006158,   0.006158,    0.006158,    0.006158,
  0.006042,   0.006042,    0.006042,    0.006042,
  0.005915,   0.005915,    0.005915,    0.005915,
  0.00584,    0.00584,     0.00584,     0.00584,
  0.005752,   0.005752,    0.005752,    0.005752,
  0.005619,   0.005619,    0.005619,    0.005619,
  0.005519,   0.005519,    0.005519,    0.005519,
  0.005451,   0.005451,    0.005451,    0.005451,
  0.005437,   0.005437,    0.005437,    0.005437,
  0.005522,   0.005522,    0.005522,    0.005522,
  0.005707,   0.005707,    0.005707,    0.005707,
  0.005897,   0.005897,    0.005897,    0.005897,
  0.006005,   0.006005,    0.006005,    0.006005,
  0.005987,   0.005987,    0.005987,    0.005987,
  0.005928,   0.005928,    0.005928,    0.005928,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005893,   0.005893,    0.005893,    0.005893,
  0.005798,   0.005798,    0.005798,    0.005798,
  0.005735,   0.005735,    0.005735,    0.005735,
  0.005784,   0.005784,    0.005784,    0.005784,
  0.005911,   0.005911,    0.005911,    0.005911,
  0.006007,   0.006007,    0.006007,    0.006007,
  0.005913,   0.005913,    0.005913,    0.005913,
  0.005783,   0.005783,    0.005783,    0.005783,
  0.005714,   0.005714,    0.005714,    0.005714,
  0.005706,   0.005706,    0.005706,    0.005706,
  0.005805,   0.005805,    0.005805,    0.005805,
  0.005951,   0.005951,    0.005951,    0.005951,
  0.006147,   0.006147,    0.006147,    0.006147,
  0.006397,   0.006397,    0.006397,    0.006397,
  0.006417,   0.006417,    0.006417,    0.006417,
  0.006121,   0.006121,    0.006121,    0.006121,
  0.006164,   0.006164,    0.006164,    0.006164,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006048,   0.006048,    0.006048,    0.006048,
  0.005859,   0.005859,    0.005859,    0.005859,
  0.005865,   0.005865,    0.005865,    0.005865,
  0.006029,   0.006029,    0.006029,    0.006029,
  0.00602,    0.00602,     0.00602,     0.00602,
  0.005988,   0.005988,    0.005988,    0.005988,
  0.006052,   0.006052,    0.006052,    0.006052,
  0.006071,   0.006071,    0.006071,    0.006071,
  0.006108,   0.006108,    0.006108,    0.006108,
  0.006126,   0.006126,    0.006126,    0.006126,
  0.006139,   0.006139,    0.006139,    0.006139,
  0.006147,   0.006147,    0.006147,    0.006147,
  0.006091,   0.006091,    0.006091,    0.006091,
  0.00606,    0.00606,     0.00606,     0.00606,
  0.006097,   0.006097,    0.006097,    0.006097,
  0.00611,    0.00611,     0.00611,     0.00611,
  0.006123,   0.006123,    0.006123,    0.006123,
  0.00611,    0.00611,     0.00611,     0.00611,
  0.00606,    0.00606,     0.00606,     0.00606,
  0.005992,   0.005992,    0.005992,    0.005992,
  0.005979,   0.005979,    0.005979,    0.005979,
  0.005979,   0.005979,    0.005979,    0.005979,
  0.005937,   0.005937,    0.005937,    0.005937,
  0.005919,   0.005919,    0.005919,    0.005919,
  0.005883,   0.005883,    0.005883,    0.005883,
  0.005773,   0.005773,    0.005773,    0.005773,
  0.005671,   0.005671,    0.005671,    0.005671,
  0.005643,   0.005643,    0.005643,    0.005643,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005486,   0.005486,    0.005486,    0.005486,
  0.005403,   0.005403,    0.005403,    0.005403,
  0.005386,   0.005386,    0.005386,    0.005386,
  0.005437,   0.005437,    0.005437,    0.005437,
  0.005505,   0.005505,    0.005505,    0.005505,
  0.005686,   0.005686,    0.005686,    0.005686,
  0.005914,   0.005914,    0.005914,    0.005914,
  0.006018,   0.006018,    0.006018,    0.006018,
  0.006016,   0.006016,    0.006016,    0.006016,
  0.005938,   0.005938,    0.005938,    0.005938,
  0.005842,   0.005842,    0.005842,    0.005842,
  0.005476,   0.005476,    0.005476,    0.005476,
  0.00504,    0.00504,     0.00504,     0.00504,
  0.004897,   0.004897,    0.004897,    0.004897,
  0.00497,    0.00497,     0.00497,     0.00497,
  0.005101,   0.005101,    0.005101,    0.005101,
  0.005491,   0.005491,    0.005491,    0.005491,
  0.005841,   0.005841,    0.005841,    0.005841,
  0.005773,   0.005773,    0.005773,    0.005773,
  0.005719,   0.005719,    0.005719,    0.005719,
  0.005784,   0.005784,    0.005784,    0.005784,
  0.005838,   0.005838,    0.005838,    0.005838,
  0.005758,   0.005758,    0.005758,    0.005758,
  0.005608,   0.005608,    0.005608,    0.005608,
  0.005586,   0.005586,    0.005586,    0.005586,
  0.005799,   0.005799,    0.005799,    0.005799,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.006102,   0.006102,    0.006102,    0.006102,
  0.006146,   0.006146,    0.006146,    0.006146,
  0.006178,   0.006178,    0.006178,    0.006178,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.006123,   0.006123,    0.006123,    0.006123,
  0.006086,   0.006086,    0.006086,    0.006086,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.006086,   0.006086,    0.006086,    0.006086,
  0.006086,   0.006086,    0.006086,    0.006086,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.006014,   0.006014,    0.006014,    0.006014,
  0.005996,   0.005996,    0.005996,    0.005996,
  0.005996,   0.005996,    0.005996,    0.005996,
  0.005996,   0.005996,    0.005996,    0.005996,
  0.005996,   0.005996,    0.005996,    0.005996,
  0.005996,   0.005996,    0.005996,    0.005996,
  0.005978,   0.005978,    0.005978,    0.005978,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.005836,   0.005836,    0.005836,    0.005836,
  0.005801,   0.005801,    0.005801,    0.005801,
  0.005766,   0.005766,    0.005766,    0.005766,
  0.005766,   0.005766,    0.005766,    0.005766,
  0.005801,   0.005801,    0.005801,    0.005801,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005906,   0.005906,    0.005906,    0.005906,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005996,   0.005996,    0.005996,    0.005996,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.00606,    0.00606,     0.00606,     0.00606,
  0.006013,   0.006013,    0.006013,    0.006013,
  0.006,      0.006,       0.006,       0.006,
  0.006071,   0.006071,    0.006071,    0.006071,
  0.006104,   0.006104,    0.006104,    0.006104,
  0.006112,   0.006112,    0.006112,    0.006112,
  0.006137,   0.006137,    0.006137,    0.006137,
  0.006079,   0.006079,    0.006079,    0.006079,
  0.006102,   0.006102,    0.006102,    0.006102,
  0.006179,   0.006179,    0.006179,    0.006179,
  0.006175,   0.006175,    0.006175,    0.006175,
  0.006184,   0.006184,    0.006184,    0.006184,
  0.006183,   0.006183,    0.006183,    0.006183,
  0.006157,   0.006157,    0.006157,    0.006157,
  0.00604,    0.00604,     0.00604,     0.00604,
  0.005863,   0.005863,    0.005863,    0.005863,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005697,   0.005697,    0.005697,    0.005697,
  0.005629,   0.005629,    0.005629,    0.005629,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005595,   0.005595,    0.005595,    0.005595,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005663,   0.005663,    0.005663,    0.005663,
  0.00568,    0.00568,     0.00568,     0.00568,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005561,   0.005561,    0.005561,    0.005561,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.00551,    0.00551,     0.00551,     0.00551,
  0.005612,   0.005612,    0.005612,    0.005612,
  0.005697,   0.005697,    0.005697,    0.005697,
  0.005714,   0.005714,    0.005714,    0.005714,
  0.005784,   0.005784,    0.005784,    0.005784,
  0.005871,   0.005871,    0.005871,    0.005871,
  0.005806,   0.005806,    0.005806,    0.005806,
  0.005603,   0.005603,    0.005603,    0.005603,
  0.005478,   0.005478,    0.005478,    0.005478,
  0.005487,   0.005487,    0.005487,    0.005487,
  0.005518,   0.005518,    0.005518,    0.005518,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.00553,    0.00553,     0.00553,     0.00553,
  0.005486,   0.005486,    0.005486,    0.005486,
  0.005433,   0.005433,    0.005433,    0.005433,
  0.005497,   0.005497,    0.005497,    0.005497,
  0.005627,   0.005627,    0.005627,    0.005627,
  0.005676,   0.005676,    0.005676,    0.005676,
  0.005676,   0.005676,    0.005676,    0.005676,
  0.005686,   0.005686,    0.005686,    0.005686,
  0.005685,   0.005685,    0.005685,    0.005685,
  0.005641,   0.005641,    0.005641,    0.005641,
  0.00568,    0.00568,     0.00568,     0.00568,
  0.00575,    0.00575,     0.00575,     0.00575,
  0.005782,   0.005782,    0.005782,    0.005782,
  0.0058,     0.0058,      0.0058,      0.0058,
  0.0058,     0.0058,      0.0058,      0.0058,
  0.005813,   0.005813,    0.005813,    0.005813,
  0.005832,   0.005832,    0.005832,    0.005832,
  0.005887,   0.005887,    0.005887,    0.005887,
  0.005943,   0.005943,    0.005943,    0.005943,
  0.005987,   0.005987,    0.005987,    0.005987,
  0.006044,   0.006044,    0.006044,    0.006044,
  0.006083,   0.006083,    0.006083,    0.006083,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.00623,    0.00623,     0.00623,     0.00623,
  0.006301,   0.006301,    0.006301,    0.006301,
  0.006392,   0.006392,    0.006392,    0.006392,
  0.006483,   0.006483,    0.006483,    0.006483,
  0.006554,   0.006554,    0.006554,    0.006554,
  0.0067,     0.0067,      0.0067,      0.0067,
  0.006792,   0.006792,    0.006792,    0.006792,
  0.006822,   0.006822,    0.006822,    0.006822,
  0.006885,   0.006885,    0.006885,    0.006885,
  0.006916,   0.006916,    0.006916,    0.006916,
  0.006957,   0.006957,    0.006957,    0.006957,
  0.00704,    0.00704,     0.00704,     0.00704,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007314,   0.007314,    0.007314,    0.007314,
  0.007487,   0.007487,    0.007487,    0.007487,
  0.0077,     0.0077,      0.0077,      0.0077,
  0.007841,   0.007841,    0.007841,    0.007841,
  0.007896,   0.007896,    0.007896,    0.007896,
  0.007937,   0.007937,    0.007937,    0.007937,
  0.008013,   0.008013,    0.008013,    0.008013,
  0.00813,    0.00813,     0.00813,     0.00813,
  0.008267,   0.008267,    0.008267,    0.008267,
  0.008372,   0.008372,    0.008372,    0.008372,
  0.008533,   0.008533,    0.008533,    0.008533,
  0.008613,   0.008613,    0.008613,    0.008613,
  0.008538,   0.008538,    0.008538,    0.008538,
  0.008486,   0.008486,    0.008486,    0.008486,
  0.008459,   0.008459,    0.008459,    0.008459,
  0.008426,   0.008426,    0.008426,    0.008426,
  0.008367,   0.008367,    0.008367,    0.008367,
  0.008339,   0.008339,    0.008339,    0.008339,
  0.008326,   0.008326,    0.008326,    0.008326,
  0.008271,   0.008271,    0.008271,    0.008271,
  0.008212,   0.008212,    0.008212,    0.008212,
  0.008147,   0.008147,    0.008147,    0.008147,
  0.008027,   0.008027,    0.008027,    0.008027,
  0.007918,   0.007918,    0.007918,    0.007918,
  0.007796,   0.007796,    0.007796,    0.007796,
  0.007677,   0.007677,    0.007677,    0.007677,
  0.007565,   0.007565,    0.007565,    0.007565,
  0.007446,   0.007446,    0.007446,    0.007446,
  0.007315,   0.007315,    0.007315,    0.007315,
  0.007239,   0.007239,    0.007239,    0.007239,
  0.007218,   0.007218,    0.007218,    0.007218,
  0.007134,   0.007134,    0.007134,    0.007134,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.006955,   0.006955,    0.006955,    0.006955,
  0.006811,   0.006811,    0.006811,    0.006811,
  0.006689,   0.006689,    0.006689,    0.006689,
  0.006601,   0.006601,    0.006601,    0.006601,
  0.006495,   0.006495,    0.006495,    0.006495,
  0.006379,   0.006379,    0.006379,    0.006379,
  0.006321,   0.006321,    0.006321,    0.006321,
  0.006264,   0.006264,    0.006264,    0.006264,
  0.006208,   0.006208,    0.006208,    0.006208,
  0.006208,   0.006208,    0.006208,    0.006208,
  0.006264,   0.006264,    0.006264,    0.006264,
  0.006335,   0.006335,    0.006335,    0.006335,
  0.006404,   0.006404,    0.006404,    0.006404,
  0.006498,   0.006498,    0.006498,    0.006498,
  0.006604,   0.006604,    0.006604,    0.006604,
  0.006721,   0.006721,    0.006721,    0.006721,
  0.006821,   0.006821,    0.006821,    0.006821,
  0.006944,   0.006944,    0.006944,    0.006944,
  0.00709,    0.00709,     0.00709,     0.00709,
  0.007185,   0.007185,    0.007185,    0.007185,
  0.007274,   0.007274,    0.007274,    0.007274,
  0.007346,   0.007346,    0.007346,    0.007346,
  0.007394,   0.007394,    0.007394,    0.007394,
  0.007415,   0.007415,    0.007415,    0.007415,
  0.007506,   0.007506,    0.007506,    0.007506,
  0.007569,   0.007569,    0.007569,    0.007569,
  0.007571,   0.007571,    0.007571,    0.007571,
  0.0077,     0.0077,      0.0077,      0.0077,
  0.007856,   0.007856,    0.007856,    0.007856,
  0.007979,   0.007979,    0.007979,    0.007979,
  0.008171,   0.008171,    0.008171,    0.008171,
  0.008351,   0.008351,    0.008351,    0.008351,
  0.008395,   0.008395,    0.008395,    0.008395,
  0.008417,   0.008417,    0.008417,    0.008417,
  0.00844,    0.00844,     0.00844,     0.00844,
  0.00843,    0.00843,     0.00843,     0.00843,
  0.008388,   0.008388,    0.008388,    0.008388,
  0.008297,   0.008297,    0.008297,    0.008297,
  0.008155,   0.008155,    0.008155,    0.008155,
  0.008074,   0.008074,    0.008074,    0.008074,
  0.008035,   0.008035,    0.008035,    0.008035,
  0.007919,   0.007919,    0.007919,    0.007919,
  0.007827,   0.007827,    0.007827,    0.007827,
  0.007813,   0.007813,    0.007813,    0.007813,
  0.007754,   0.007754,    0.007754,    0.007754,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007531,   0.007531,    0.007531,    0.007531,
  0.007465,   0.007465,    0.007465,    0.007465,
  0.0074,     0.0074,      0.0074,      0.0074,
  0.007421,   0.007421,    0.007421,    0.007421,
  0.007421,   0.007421,    0.007421,    0.007421,
  0.007292,   0.007292,    0.007292,    0.007292,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.007019,   0.007019,    0.007019,    0.007019,
  0.006978,   0.006978,    0.006978,    0.006978,
  0.006937,   0.006937,    0.006937,    0.006937,
  0.006896,   0.006896,    0.006896,    0.006896,
  0.006835,   0.006835,    0.006835,    0.006835,
  0.006795,   0.006795,    0.006795,    0.006795,
  0.006876,   0.006876,    0.006876,    0.006876,
  0.007125,   0.007125,    0.007125,    0.007125,
  0.007502,   0.007502,    0.007502,    0.007502,
  0.007835,   0.007835,    0.007835,    0.007835,
  0.008047,   0.008047,    0.008047,    0.008047,
  0.008176,   0.008176,    0.008176,    0.008176,
  0.008209,   0.008209,    0.008209,    0.008209,
  0.008257,   0.008257,    0.008257,    0.008257,
  0.008349,   0.008349,    0.008349,    0.008349,
  0.008409,   0.008409,    0.008409,    0.008409,
  0.008489,   0.008489,    0.008489,    0.008489,
  0.008547,   0.008547,    0.008547,    0.008547,
  0.008455,   0.008455,    0.008455,    0.008455,
  0.008392,   0.008392,    0.008392,    0.008392,
  0.008519,   0.008519,    0.008519,    0.008519,
  0.008647,   0.008647,    0.008647,    0.008647,
  0.008738,   0.008738,    0.008738,    0.008738,
  0.008892,   0.008892,    0.008892,    0.008892,
  0.00896,    0.00896,     0.00896,     0.00896,
  0.008905,   0.008905,    0.008905,    0.008905,
  0.008902,   0.008902,    0.008902,    0.008902,
  0.008973,   0.008973,    0.008973,    0.008973,
  0.009101,   0.009101,    0.009101,    0.009101,
  0.009092,   0.009092,    0.009092,    0.009092,
  0.008897,   0.008897,    0.008897,    0.008897,
  0.008666,   0.008666,    0.008666,    0.008666,
  0.00839,    0.00839,     0.00839,     0.00839,
  0.008146,   0.008146,    0.008146,    0.008146,
  0.007914,   0.007914,    0.007914,    0.007914,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007296,   0.007296,    0.007296,    0.007296,
  0.006917,   0.006917,    0.006917,    0.006917,
  0.007022,   0.007022,    0.007022,    0.007022,
  0.007423,   0.007423,    0.007423,    0.007423,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007777,   0.007777,    0.007777,    0.007777,
  0.007982,   0.007982,    0.007982,    0.007982,
  0.008075,   0.008075,    0.008075,    0.008075,
  0.008075,   0.008075,    0.008075,    0.008075,
  0.008028,   0.008028,    0.008028,    0.008028,
  0.008005,   0.008005,    0.008005,    0.008005,
  0.007982,   0.007982,    0.007982,    0.007982,
  0.007959,   0.007959,    0.007959,    0.007959,
  0.007959,   0.007959,    0.007959,    0.007959,
  0.00777,    0.00777,     0.00777,     0.00777,
  0.007449,   0.007449,    0.007449,    0.007449,
  0.007295,   0.007295,    0.007295,    0.007295,
  0.007249,   0.007249,    0.007249,    0.007249,
  0.007062,   0.007062,    0.007062,    0.007062,
  0.006654,   0.006654,    0.006654,    0.006654,
  0.006242,   0.006242,    0.006242,    0.006242,
  0.005842,   0.005842,    0.005842,    0.005842,
  0.005516,   0.005516,    0.005516,    0.005516,
  0.00538,    0.00538,     0.00538,     0.00538,
  0.005286,   0.005286,    0.005286,    0.005286,
  0.005223,   0.005223,    0.005223,    0.005223,
  0.005202,   0.005202,    0.005202,    0.005202,
  0.005159,   0.005159,    0.005159,    0.005159,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.004761,   0.004761,    0.004761,    0.004761,
  0.004488,   0.004488,    0.004488,    0.004488,
  0.004257,   0.004257,    0.004257,    0.004257,
  0.004141,   0.004141,    0.004141,    0.004141,
  0.004184,   0.004184,    0.004184,    0.004184,
  0.004281,   0.004281,    0.004281,    0.004281,
  0.00431,    0.00431,     0.00431,     0.00431,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004353,   0.004353,    0.004353,    0.004353,
  0.00444,    0.00444,     0.00444,     0.00444,
  0.004466,   0.004466,    0.004466,    0.004466,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.00448,    0.00448,     0.00448,     0.00448,
  0.004446,   0.004446,    0.004446,    0.004446,
  0.004399,   0.004399,    0.004399,    0.004399,
  0.004399,   0.004399,    0.004399,    0.004399,
  0.004414,   0.004414,    0.004414,    0.004414,
  0.00435,    0.00435,     0.00435,     0.00435,
  0.004271,   0.004271,    0.004271,    0.004271,
  0.00424,    0.00424,     0.00424,     0.00424,
  0.004225,   0.004225,    0.004225,    0.004225,
  0.004227,   0.004227,    0.004227,    0.004227,
  0.004199,   0.004199,    0.004199,    0.004199,
  0.004126,   0.004126,    0.004126,    0.004126,
  0.004073,   0.004073,    0.004073,    0.004073,
  0.004018,   0.004018,    0.004018,    0.004018,
  0.003961,   0.003961,    0.003961,    0.003961,
  0.003902,   0.003902,    0.003902,    0.003902,
  0.003853,   0.003853,    0.003853,    0.003853,
  0.003811,   0.003811,    0.003811,    0.003811,
  0.003778,   0.003778,    0.003778,    0.003778,
  0.003728,   0.003728,    0.003728,    0.003728,
  0.00368,    0.00368,     0.00368,     0.00368,
  0.003659,   0.003659,    0.003659,    0.003659,
  0.003646,   0.003646,    0.003646,    0.003646,
  0.003659,   0.003659,    0.003659,    0.003659,
  0.003685,   0.003685,    0.003685,    0.003685,
  0.003711,   0.003711,    0.003711,    0.003711,
  0.003778,   0.003778,    0.003778,    0.003778,
  0.003856,   0.003856,    0.003856,    0.003856,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003978,   0.003978,    0.003978,    0.003978,
  0.003994,   0.003994,    0.003994,    0.003994,
  0.003974,   0.003974,    0.003974,    0.003974,
  0.003927,   0.003927,    0.003927,    0.003927,
  0.003816,   0.003816,    0.003816,    0.003816,
  0.003637,   0.003637,    0.003637,    0.003637,
  0.003531,   0.003531,    0.003531,    0.003531,
  0.00347,    0.00347,     0.00347,     0.00347,
  0.003434,   0.003434,    0.003434,    0.003434,
  0.003431,   0.003431,    0.003431,    0.003431,
  0.003462,   0.003462,    0.003462,    0.003462,
  0.00356,    0.00356,     0.00356,     0.00356,
  0.003652,   0.003652,    0.003652,    0.003652,
  0.003751,   0.003751,    0.003751,    0.003751,
  0.003938,   0.003938,    0.003938,    0.003938,
  0.004108,   0.004108,    0.004108,    0.004108,
  0.00421,    0.00421,     0.00421,     0.00421,
  0.004244,   0.004244,    0.004244,    0.004244,
  0.004194,   0.004194,    0.004194,    0.004194,
  0.004104,   0.004104,    0.004104,    0.004104,
  0.004005,   0.004005,    0.004005,    0.004005,
  0.003932,   0.003932,    0.003932,    0.003932,
  0.003918,   0.003918,    0.003918,    0.003918,
  0.003892,   0.003892,    0.003892,    0.003892,
  0.003835,   0.003835,    0.003835,    0.003835,
  0.003755,   0.003755,    0.003755,    0.003755,
  0.003675,   0.003675,    0.003675,    0.003675,
  0.003605,   0.003605,    0.003605,    0.003605,
  0.003558,   0.003558,    0.003558,    0.003558,
  0.003549,   0.003549,    0.003549,    0.003549,
  0.003513,   0.003513,    0.003513,    0.003513,
  0.003481,   0.003481,    0.003481,    0.003481,
  0.003499,   0.003499,    0.003499,    0.003499,
  0.003494,   0.003494,    0.003494,    0.003494,
  0.003485,   0.003485,    0.003485,    0.003485,
  0.003488,   0.003488,    0.003488,    0.003488,
  0.003464,   0.003464,    0.003464,    0.003464,
  0.003433,   0.003433,    0.003433,    0.003433,
  0.003433,   0.003433,    0.003433,    0.003433,
  0.003445,   0.003445,    0.003445,    0.003445,
  0.003418,   0.003418,    0.003418,    0.003418,
  0.003391,   0.003391,    0.003391,    0.003391,
  0.003374,   0.003374,    0.003374,    0.003374,
  0.003354,   0.003354,    0.003354,    0.003354,
  0.003366,   0.003366,    0.003366,    0.003366,
  0.003442,   0.003442,    0.003442,    0.003442,
  0.003553,   0.003553,    0.003553,    0.003553,
  0.003631,   0.003631,    0.003631,    0.003631,
  0.003646,   0.003646,    0.003646,    0.003646,
  0.003618,   0.003618,    0.003618,    0.003618,
  0.003581,   0.003581,    0.003581,    0.003581,
  0.003584,   0.003584,    0.003584,    0.003584,
  0.00363,    0.00363,     0.00363,     0.00363,
  0.003538,   0.003538,    0.003538,    0.003538,
  0.003318,   0.003318,    0.003318,    0.003318,
  0.003222,   0.003222,    0.003222,    0.003222,
  0.003141,   0.003141,    0.003141,    0.003141,
  0.003126,   0.003126,    0.003126,    0.003126,
  0.003196,   0.003196,    0.003196,    0.003196,
  0.003175,   0.003175,    0.003175,    0.003175,
  0.003302,   0.003302,    0.003302,    0.003302,
  0.003551,   0.003551,    0.003551,    0.003551,
  0.003705,   0.003705,    0.003705,    0.003705,
  0.003759,   0.003759,    0.003759,    0.003759,
  0.003744,   0.003744,    0.003744,    0.003744,
  0.003726,   0.003726,    0.003726,    0.003726,
  0.003764,   0.003764,    0.003764,    0.003764,
  0.003883,   0.003883,    0.003883,    0.003883,
  0.003988,   0.003988,    0.003988,    0.003988,
  0.004075,   0.004075,    0.004075,    0.004075,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.004063,   0.004063,    0.004063,    0.004063,
  0.00408,    0.00408,     0.00408,     0.00408,
  0.004106,   0.004106,    0.004106,    0.004106,
  0.00403,    0.00403,     0.00403,     0.00403,
  0.004039,   0.004039,    0.004039,    0.004039,
  0.00413,    0.00413,     0.00413,     0.00413,
  0.004108,   0.004108,    0.004108,    0.004108,
  0.004102,   0.004102,    0.004102,    0.004102,
  0.004095,   0.004095,    0.004095,    0.004095,
  0.004081,   0.004081,    0.004081,    0.004081,
  0.004042,   0.004042,    0.004042,    0.004042,
  0.004074,   0.004074,    0.004074,    0.004074,
  0.00417,    0.00417,     0.00417,     0.00417,
  0.004181,   0.004181,    0.004181,    0.004181,
  0.004196,   0.004196,    0.004196,    0.004196,
  0.004196,   0.004196,    0.004196,    0.004196,
  0.004187,   0.004187,    0.004187,    0.004187,
  0.004247,   0.004247,    0.004247,    0.004247,
  0.004317,   0.004317,    0.004317,    0.004317,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004436,   0.004436,    0.004436,    0.004436,
  0.004512,   0.004512,    0.004512,    0.004512,
  0.004652,   0.004652,    0.004652,    0.004652,
  0.004855,   0.004855,    0.004855,    0.004855,
  0.005097,   0.005097,    0.005097,    0.005097,
  0.005437,   0.005437,    0.005437,    0.005437,
  0.005784,   0.005784,    0.005784,    0.005784,
  0.00595,    0.00595,     0.00595,     0.00595,
  0.00572,    0.00572,     0.00572,     0.00572,
  0.005244,   0.005244,    0.005244,    0.005244,
  0.004929,   0.004929,    0.004929,    0.004929,
  0.004876,   0.004876,    0.004876,    0.004876,
  0.004981,   0.004981,    0.004981,    0.004981,
  0.005033,   0.005033,    0.005033,    0.005033,
  0.005033,   0.005033,    0.005033,    0.005033,
  0.005076,   0.005076,    0.005076,    0.005076,
  0.005128,   0.005128,    0.005128,    0.005128,
  0.005193,   0.005193,    0.005193,    0.005193,
  0.005295,   0.005295,    0.005295,    0.005295,
  0.005361,   0.005361,    0.005361,    0.005361,
  0.00537,    0.00537,     0.00537,     0.00537,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005461,   0.005461,    0.005461,    0.005461,
  0.005524,   0.005524,    0.005524,    0.005524,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.00565,    0.00565,     0.00565,     0.00565,
  0.005647,   0.005647,    0.005647,    0.005647,
  0.005612,   0.005612,    0.005612,    0.005612,
  0.005557,   0.005557,    0.005557,    0.005557,
  0.005519,   0.005519,    0.005519,    0.005519,
  0.005502,   0.005502,    0.005502,    0.005502,
  0.005483,   0.005483,    0.005483,    0.005483,
  0.005512,   0.005512,    0.005512,    0.005512,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005648,   0.005648,    0.005648,    0.005648,
  0.005571,   0.005571,    0.005571,    0.005571,
  0.005408,   0.005408,    0.005408,    0.005408,
  0.005257,   0.005257,    0.005257,    0.005257,
  0.005077,   0.005077,    0.005077,    0.005077,
  0.004871,   0.004871,    0.004871,    0.004871,
  0.00476,    0.00476,     0.00476,     0.00476,
  0.004681,   0.004681,    0.004681,    0.004681,
  0.004527,   0.004527,    0.004527,    0.004527,
  0.004391,   0.004391,    0.004391,    0.004391,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004354,   0.004354,    0.004354,    0.004354,
  0.004291,   0.004291,    0.004291,    0.004291,
  0.004298,   0.004298,    0.004298,    0.004298,
  0.004379,   0.004379,    0.004379,    0.004379,
  0.004536,   0.004536,    0.004536,    0.004536,
  0.004825,   0.004825,    0.004825,    0.004825,
  0.00508,    0.00508,     0.00508,     0.00508,
  0.005198,   0.005198,    0.005198,    0.005198,
  0.005291,   0.005291,    0.005291,    0.005291,
  0.005196,   0.005196,    0.005196,    0.005196,
  0.004904,   0.004904,    0.004904,    0.004904,
  0.004658,   0.004658,    0.004658,    0.004658,
  0.004515,   0.004515,    0.004515,    0.004515,
  0.004435,   0.004435,    0.004435,    0.004435,
  0.004356,   0.004356,    0.004356,    0.004356,
  0.004066,   0.004066,    0.004066,    0.004066,
  0.003825,   0.003825,    0.003825,    0.003825,
  0.003939,   0.003939,    0.003939,    0.003939,
  0.004132,   0.004132,    0.004132,    0.004132,
  0.004314,   0.004314,    0.004314,    0.004314,
  0.004419,   0.004419,    0.004419,    0.004419,
  0.004439,   0.004439,    0.004439,    0.004439,
  0.004475,   0.004475,    0.004475,    0.004475,
  0.004548,   0.004548,    0.004548,    0.004548,
  0.004595,   0.004595,    0.004595,    0.004595,
  0.004647,   0.004647,    0.004647,    0.004647,
  0.004721,   0.004721,    0.004721,    0.004721,
  0.004766,   0.004766,    0.004766,    0.004766,
  0.004826,   0.004826,    0.004826,    0.004826,
  0.004871,   0.004871,    0.004871,    0.004871,
  0.00487,    0.00487,     0.00487,     0.00487,
  0.004901,   0.004901,    0.004901,    0.004901,
  0.004901,   0.004901,    0.004901,    0.004901,
  0.004886,   0.004886,    0.004886,    0.004886,
  0.004918,   0.004918,    0.004918,    0.004918,
  0.004933,   0.004933,    0.004933,    0.004933,
  0.004949,   0.004949,    0.004949,    0.004949,
  0.004919,   0.004919,    0.004919,    0.004919,
  0.004846,   0.004846,    0.004846,    0.004846,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004788,   0.004788,    0.004788,    0.004788,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004671,   0.004671,    0.004671,    0.004671,
  0.004656,   0.004656,    0.004656,    0.004656,
  0.004671,   0.004671,    0.004671,    0.004671,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005395,   0.005395,    0.005395,    0.005395,
  0.005547,   0.005547,    0.005547,    0.005547,
  0.005637,   0.005637,    0.005637,    0.005637,
  0.005687,   0.005687,    0.005687,    0.005687,
  0.005722,   0.005722,    0.005722,    0.005722,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005713,   0.005713,    0.005713,    0.005713,
  0.005639,   0.005639,    0.005639,    0.005639,
  0.005553,   0.005553,    0.005553,    0.005553,
  0.005418,   0.005418,    0.005418,    0.005418,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005275,   0.005275,    0.005275,    0.005275,
  0.005307,   0.005307,    0.005307,    0.005307,
  0.005433,   0.005433,    0.005433,    0.005433,
  0.00559,    0.00559,     0.00559,     0.00559,
  0.005674,   0.005674,    0.005674,    0.005674,
  0.005717,   0.005717,    0.005717,    0.005717,
  0.005943,   0.005943,    0.005943,    0.005943,
  0.006212,   0.006212,    0.006212,    0.006212,
  0.006283,   0.006283,    0.006283,    0.006283,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006234,   0.006234,    0.006234,    0.006234,
  0.006215,   0.006215,    0.006215,    0.006215,
  0.006197,   0.006197,    0.006197,    0.006197,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.005978,   0.005978,    0.005978,    0.005978,
  0.005928,   0.005928,    0.005928,    0.005928,
  0.005847,   0.005847,    0.005847,    0.005847,
  0.005704,   0.005704,    0.005704,    0.005704,
  0.005546,   0.005546,    0.005546,    0.005546,
  0.00542,    0.00542,     0.00542,     0.00542,
  0.005326,   0.005326,    0.005326,    0.005326,
  0.005395,   0.005395,    0.005395,    0.005395,
  0.005525,   0.005525,    0.005525,    0.005525,
  0.005551,   0.005551,    0.005551,    0.005551,
  0.005563,   0.005563,    0.005563,    0.005563,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.005444,   0.005444,    0.005444,    0.005444,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005394,   0.005394,    0.005394,    0.005394,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.00556,    0.00556,     0.00556,     0.00556,
  0.005646,   0.005646,    0.005646,    0.005646,
  0.005855,   0.005855,    0.005855,    0.005855,
  0.006105,   0.006105,    0.006105,    0.006105,
  0.006241,   0.006241,    0.006241,    0.006241,
  0.006164,   0.006164,    0.006164,    0.006164,
  0.005985,   0.005985,    0.005985,    0.005985,
  0.005812,   0.005812,    0.005812,    0.005812,
  0.005695,   0.005695,    0.005695,    0.005695,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005455,   0.005455,    0.005455,    0.005455,
  0.005455,   0.005455,    0.005455,    0.005455,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005854,   0.005854,    0.005854,    0.005854,
  0.006034,   0.006034,    0.006034,    0.006034,
  0.006059,   0.006059,    0.006059,    0.006059,
  0.006128,   0.006128,    0.006128,    0.006128,
  0.006163,   0.006163,    0.006163,    0.006163,
  0.006179,   0.006179,    0.006179,    0.006179,
  0.006196,   0.006196,    0.006196,    0.006196,
  0.006202,   0.006202,    0.006202,    0.006202,
  0.00622,    0.00622,     0.00622,     0.00622,
  0.006239,   0.006239,    0.006239,    0.006239,
  0.006234,   0.006234,    0.006234,    0.006234,
  0.006197,   0.006197,    0.006197,    0.006197,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.006105,   0.006105,    0.006105,    0.006105,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.005818,   0.005818,    0.005818,    0.005818,
  0.005748,   0.005748,    0.005748,    0.005748,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005444,   0.005444,    0.005444,    0.005444,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005249,   0.005249,    0.005249,    0.005249,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.004918,   0.004918,    0.004918,    0.004918,
  0.004704,   0.004704,    0.004704,    0.004704,
  0.004452,   0.004452,    0.004452,    0.004452,
  0.004158,   0.004158,    0.004158,    0.004158,
  0.003931,   0.003931,    0.003931,    0.003931,
  0.003843,   0.003843,    0.003843,    0.003843,
  0.003752,   0.003752,    0.003752,    0.003752,
  0.003631,   0.003631,    0.003631,    0.003631,
  0.003555,   0.003555,    0.003555,    0.003555,
  0.003506,   0.003506,    0.003506,    0.003506,
  0.00346,    0.00346,     0.00346,     0.00346,
  0.003351,   0.003351,    0.003351,    0.003351,
  0.003249,   0.003249,    0.003249,    0.003249,
  0.003136,   0.003136,    0.003136,    0.003136,
  0.00289,    0.00289,     0.00289,     0.00289,
  0.00265,    0.00265,     0.00265,     0.00265,
  0.002539,   0.002539,    0.002539,    0.002539,
  0.002476,   0.002476,    0.002476,    0.002476,
  0.00243,    0.00243,     0.00243,     0.00243,
  0.0024,     0.0024,      0.0024,      0.0024,
  0.002449,   0.002449,    0.002449,    0.002449,
  0.002481,   0.002481,    0.002481,    0.002481,
  0.002402,   0.002402,    0.002402,    0.002402,
  0.002322,   0.002322,    0.002322,    0.002322,
  0.002321,   0.002321,    0.002321,    0.002321,
  0.002398,   0.002398,    0.002398,    0.002398,
  0.00251,    0.00251,     0.00251,     0.00251,
  0.002601,   0.002601,    0.002601,    0.002601,
  0.00265,    0.00265,     0.00265,     0.00265,
  0.002646,   0.002646,    0.002646,    0.002646,
  0.002712,   0.002712,    0.002712,    0.002712,
  0.002942,   0.002942,    0.002942,    0.002942,
  0.003084,   0.003084,    0.003084,    0.003084,
  0.003065,   0.003065,    0.003065,    0.003065,
  0.003045,   0.003045,    0.003045,    0.003045,
  0.003058,   0.003058,    0.003058,    0.003058,
  0.00309,    0.00309,     0.00309,     0.00309,
  0.003111,   0.003111,    0.003111,    0.003111,
  0.003071,   0.003071,    0.003071,    0.003071,
  0.00302,    0.00302,     0.00302,     0.00302,
  0.003024,   0.003024,    0.003024,    0.003024,
  0.003021,   0.003021,    0.003021,    0.003021,
  0.002976,   0.002976,    0.002976,    0.002976,
  0.002951,   0.002951,    0.002951,    0.002951,
  0.002938,   0.002938,    0.002938,    0.002938,
  0.002907,   0.002907,    0.002907,    0.002907,
  0.002898,   0.002898,    0.002898,    0.002898,
  0.002898,   0.002898,    0.002898,    0.002898,
  0.002886,   0.002886,    0.002886,    0.002886,
  0.002864,   0.002864,    0.002864,    0.002864,
  0.002832,   0.002832,    0.002832,    0.002832,
  0.002821,   0.002821,    0.002821,    0.002821,
  0.002821,   0.002821,    0.002821,    0.002821,
  0.00281,    0.00281,     0.00281,     0.00281,
  0.00281,    0.00281,     0.00281,     0.00281,
  0.002799,   0.002799,    0.002799,    0.002799,
  0.00281,    0.00281,     0.00281,     0.00281,
  0.00286,    0.00286,     0.00286,     0.00286,
  0.002889,   0.002889,    0.002889,    0.002889,
  0.002864,   0.002864,    0.002864,    0.002864,
  0.002835,   0.002835,    0.002835,    0.002835,
  0.002809,   0.002809,    0.002809,    0.002809,
  0.002757,   0.002757,    0.002757,    0.002757,
  0.002798,   0.002798,    0.002798,    0.002798,
  0.002714,   0.002714,    0.002714,    0.002714,
  0.002555,   0.002555,    0.002555,    0.002555,
  0.002508,   0.002508,    0.002508,    0.002508,
  0.002415,   0.002415,    0.002415,    0.002415,
  0.002339,   0.002339,    0.002339,    0.002339,
  0.002325,   0.002325,    0.002325,    0.002325,
  0.002327,   0.002327,    0.002327,    0.002327,
  0.002295,   0.002295,    0.002295,    0.002295,
  0.002309,   0.002309,    0.002309,    0.002309,
  0.002431,   0.002431,    0.002431,    0.002431,
  0.002638,   0.002638,    0.002638,    0.002638,
  0.00278,    0.00278,     0.00278,     0.00278,
  0.002727,   0.002727,    0.002727,    0.002727,
  0.002648,   0.002648,    0.002648,    0.002648,
  0.002634,   0.002634,    0.002634,    0.002634,
  0.002631,   0.002631,    0.002631,    0.002631,
  0.002676,   0.002676,    0.002676,    0.002676,
  0.002731,   0.002731,    0.002731,    0.002731,
  0.002731,   0.002731,    0.002731,    0.002731,
  0.002744,   0.002744,    0.002744,    0.002744,
  0.002751,   0.002751,    0.002751,    0.002751,
  0.002729,   0.002729,    0.002729,    0.002729,
  0.002748,   0.002748,    0.002748,    0.002748,
  0.002761,   0.002761,    0.002761,    0.002761,
  0.002747,   0.002747,    0.002747,    0.002747,
  0.002726,   0.002726,    0.002726,    0.002726,
  0.002706,   0.002706,    0.002706,    0.002706,
  0.002702,   0.002702,    0.002702,    0.002702,
  0.002717,   0.002717,    0.002717,    0.002717,
  0.002746,   0.002746,    0.002746,    0.002746,
  0.002735,   0.002735,    0.002735,    0.002735,
  0.002725,   0.002725,    0.002725,    0.002725,
  0.002735,   0.002735,    0.002735,    0.002735,
  0.002703,   0.002703,    0.002703,    0.002703,
  0.002662,   0.002662,    0.002662,    0.002662,
  0.002642,   0.002642,    0.002642,    0.002642,
  0.00261,    0.00261,     0.00261,     0.00261,
  0.002589,   0.002589,    0.002589,    0.002589,
  0.002602,   0.002602,    0.002602,    0.002602,
  0.002612,   0.002612,    0.002612,    0.002612,
  0.002588,   0.002588,    0.002588,    0.002588,
  0.002599,   0.002599,    0.002599,    0.002599,
  0.002668,   0.002668,    0.002668,    0.002668,
  0.002714,   0.002714,    0.002714,    0.002714,
  0.002756,   0.002756,    0.002756,    0.002756,
  0.002763,   0.002763,    0.002763,    0.002763,
  0.00267,    0.00267,     0.00267,     0.00267,
  0.002495,   0.002495,    0.002495,    0.002495,
  0.002264,   0.002264,    0.002264,    0.002264,
  0.002069,   0.002069,    0.002069,    0.002069,
  0.001962,   0.001962,    0.001962,    0.001962,
  0.001869,   0.001869,    0.001869,    0.001869,
  0.001645,   0.001645,    0.001645,    0.001645,
  0.001485,   0.001485,    0.001485,    0.001485,
  0.001574,   0.001574,    0.001574,    0.001574,
  0.001608,   0.001608,    0.001608,    0.001608,
  0.002041,   0.002041,    0.002041,    0.002041,
  0.002626,   0.002626,    0.002626,    0.002626,
  0.002746,   0.002746,    0.002746,    0.002746,
  0.002784,   0.002784,    0.002784,    0.002784,
  0.002793,   0.002793,    0.002793,    0.002793,
  0.002784,   0.002784,    0.002784,    0.002784,
  0.002752,   0.002752,    0.002752,    0.002752,
  0.002738,   0.002738,    0.002738,    0.002738,
  0.002712,   0.002712,    0.002712,    0.002712,
  0.002624,   0.002624,    0.002624,    0.002624,
  0.002559,   0.002559,    0.002559,    0.002559,
  0.002535,   0.002535,    0.002535,    0.002535,
  0.00256,    0.00256,     0.00256,     0.00256,
  0.002566,   0.002566,    0.002566,    0.002566,
  0.002561,   0.002561,    0.002561,    0.002561,
  0.002555,   0.002555,    0.002555,    0.002555,
  0.002435,   0.002435,    0.002435,    0.002435,
  0.002265,   0.002265,    0.002265,    0.002265,
  0.002253,   0.002253,    0.002253,    0.002253,
  0.002359,   0.002359,    0.002359,    0.002359,
  0.002434,   0.002434,    0.002434,    0.002434,
  0.002485,   0.002485,    0.002485,    0.002485,
  0.002504,   0.002504,    0.002504,    0.002504,
  0.002478,   0.002478,    0.002478,    0.002478,
  0.002466,   0.002466,    0.002466,    0.002466,
  0.002435,   0.002435,    0.002435,    0.002435,
  0.002485,   0.002485,    0.002485,    0.002485,
  0.002586,   0.002586,    0.002586,    0.002586,
  0.002644,   0.002644,    0.002644,    0.002644,
  0.002739,   0.002739,    0.002739,    0.002739,
  0.002819,   0.002819,    0.002819,    0.002819,
  0.002869,   0.002869,    0.002869,    0.002869,
  0.002869,   0.002869,    0.002869,    0.002869,
  0.002876,   0.002876,    0.002876,    0.002876,
  0.00293,    0.00293,     0.00293,     0.00293,
  0.002974,   0.002974,    0.002974,    0.002974,
  0.00304,    0.00304,     0.00304,     0.00304,
  0.003098,   0.003098,    0.003098,    0.003098,
  0.003065,   0.003065,    0.003065,    0.003065,
  0.002921,   0.002921,    0.002921,    0.002921,
  0.002621,   0.002621,    0.002621,    0.002621,
  0.002411,   0.002411,    0.002411,    0.002411,
  0.002461,   0.002461,    0.002461,    0.002461,
  0.002597,   0.002597,    0.002597,    0.002597,
  0.002747,   0.002747,    0.002747,    0.002747,
  0.002874,   0.002874,    0.002874,    0.002874,
  0.003029,   0.003029,    0.003029,    0.003029,
  0.003049,   0.003049,    0.003049,    0.003049,
  0.003022,   0.003022,    0.003022,    0.003022,
  0.003223,   0.003223,    0.003223,    0.003223,
  0.003427,   0.003427,    0.003427,    0.003427,
  0.003497,   0.003497,    0.003497,    0.003497,
  0.003468,   0.003468,    0.003468,    0.003468,
  0.003393,   0.003393,    0.003393,    0.003393,
  0.003358,   0.003358,    0.003358,    0.003358,
  0.00339,    0.00339,     0.00339,     0.00339,
  0.003453,   0.003453,    0.003453,    0.003453,
  0.0035,     0.0035,      0.0035,      0.0035,
  0.003579,   0.003579,    0.003579,    0.003579,
  0.003675,   0.003675,    0.003675,    0.003675,
  0.003722,   0.003722,    0.003722,    0.003722,
  0.003767,   0.003767,    0.003767,    0.003767,
  0.003799,   0.003799,    0.003799,    0.003799,
  0.0038,     0.0038,      0.0038,      0.0038,
  0.003785,   0.003785,    0.003785,    0.003785,
  0.003771,   0.003771,    0.003771,    0.003771,
  0.003774,   0.003774,    0.003774,    0.003774,
  0.003751,   0.003751,    0.003751,    0.003751,
  0.003721,   0.003721,    0.003721,    0.003721,
  0.003744,   0.003744,    0.003744,    0.003744,
  0.00379,    0.00379,     0.00379,     0.00379,
  0.00378,    0.00378,     0.00378,     0.00378,
  0.00376,    0.00376,     0.00376,     0.00376,
  0.003687,   0.003687,    0.003687,    0.003687,
  0.003633,   0.003633,    0.003633,    0.003633,
  0.003671,   0.003671,    0.003671,    0.003671,
  0.003804,   0.003804,    0.003804,    0.003804,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.004012,   0.004012,    0.004012,    0.004012,
  0.004108,   0.004108,    0.004108,    0.004108,
  0.004191,   0.004191,    0.004191,    0.004191,
  0.004205,   0.004205,    0.004205,    0.004205,
  0.004195,   0.004195,    0.004195,    0.004195,
  0.00418,    0.00418,     0.00418,     0.00418,
  0.004207,   0.004207,    0.004207,    0.004207,
  0.004168,   0.004168,    0.004168,    0.004168,
  0.004121,   0.004121,    0.004121,    0.004121,
  0.004142,   0.004142,    0.004142,    0.004142,
  0.00416,    0.00416,     0.00416,     0.00416,
  0.004188,   0.004188,    0.004188,    0.004188,
  0.004173,   0.004173,    0.004173,    0.004173,
  0.004081,   0.004081,    0.004081,    0.004081,
  0.003978,   0.003978,    0.003978,    0.003978,
  0.003937,   0.003937,    0.003937,    0.003937,
  0.003978,   0.003978,    0.003978,    0.003978,
  0.003986,   0.003986,    0.003986,    0.003986,
  0.003931,   0.003931,    0.003931,    0.003931,
  0.003944,   0.003944,    0.003944,    0.003944,
  0.004051,   0.004051,    0.004051,    0.004051,
  0.004219,   0.004219,    0.004219,    0.004219,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004395,   0.004395,    0.004395,    0.004395,
  0.004424,   0.004424,    0.004424,    0.004424,
  0.004488,   0.004488,    0.004488,    0.004488,
  0.004532,   0.004532,    0.004532,    0.004532,
  0.004544,   0.004544,    0.004544,    0.004544,
  0.00454,    0.00454,     0.00454,     0.00454,
  0.004515,   0.004515,    0.004515,    0.004515,
  0.004511,   0.004511,    0.004511,    0.004511,
  0.004502,   0.004502,    0.004502,    0.004502,
  0.004462,   0.004462,    0.004462,    0.004462,
  0.0044,     0.0044,      0.0044,      0.0044,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004309,   0.004309,    0.004309,    0.004309,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004309,   0.004309,    0.004309,    0.004309,
  0.004317,   0.004317,    0.004317,    0.004317,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004291,   0.004291,    0.004291,    0.004291,
  0.004246,   0.004246,    0.004246,    0.004246,
  0.004201,   0.004201,    0.004201,    0.004201,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004238,   0.004238,    0.004238,    0.004238,
  0.004248,   0.004248,    0.004248,    0.004248,
  0.004273,   0.004273,    0.004273,    0.004273,
  0.004284,   0.004284,    0.004284,    0.004284,
  0.004267,   0.004267,    0.004267,    0.004267,
  0.00425,    0.00425,     0.00425,     0.00425,
  0.004232,   0.004232,    0.004232,    0.004232,
  0.004196,   0.004196,    0.004196,    0.004196,
  0.004191,   0.004191,    0.004191,    0.004191,
  0.004187,   0.004187,    0.004187,    0.004187,
  0.004182,   0.004182,    0.004182,    0.004182,
  0.004199,   0.004199,    0.004199,    0.004199,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004191,   0.004191,    0.004191,    0.004191,
  0.004149,   0.004149,    0.004149,    0.004149,
  0.004058,   0.004058,    0.004058,    0.004058,
  0.004024,   0.004024,    0.004024,    0.004024,
  0.003947,   0.003947,    0.003947,    0.003947,
  0.003817,   0.003817,    0.003817,    0.003817,
  0.003752,   0.003752,    0.003752,    0.003752,
  0.003693,   0.003693,    0.003693,    0.003693,
  0.0036,     0.0036,      0.0036,      0.0036,
  0.003509,   0.003509,    0.003509,    0.003509,
  0.003476,   0.003476,    0.003476,    0.003476,
  0.003443,   0.003443,    0.003443,    0.003443,
  0.003356,   0.003356,    0.003356,    0.003356,
  0.003239,   0.003239,    0.003239,    0.003239,
  0.003146,   0.003146,    0.003146,    0.003146,
  0.003095,   0.003095,    0.003095,    0.003095,
  0.003085,   0.003085,    0.003085,    0.003085,
  0.003126,   0.003126,    0.003126,    0.003126,
  0.003187,   0.003187,    0.003187,    0.003187,
  0.003249,   0.003249,    0.003249,    0.003249,
  0.003302,   0.003302,    0.003302,    0.003302,
  0.003399,   0.003399,    0.003399,    0.003399,
  0.003498,   0.003498,    0.003498,    0.003498,
  0.003532,   0.003532,    0.003532,    0.003532,
  0.003554,   0.003554,    0.003554,    0.003554,
  0.003566,   0.003566,    0.003566,    0.003566,
  0.003566,   0.003566,    0.003566,    0.003566,
  0.003577,   0.003577,    0.003577,    0.003577,
  0.003588,   0.003588,    0.003588,    0.003588,
  0.003577,   0.003577,    0.003577,    0.003577,
  0.003554,   0.003554,    0.003554,    0.003554,
  0.003543,   0.003543,    0.003543,    0.003543,
  0.003554,   0.003554,    0.003554,    0.003554,
  0.003532,   0.003532,    0.003532,    0.003532,
  0.003509,   0.003509,    0.003509,    0.003509,
  0.003566,   0.003566,    0.003566,    0.003566,
  0.003646,   0.003646,    0.003646,    0.003646,
  0.003728,   0.003728,    0.003728,    0.003728,
  0.003873,   0.003873,    0.003873,    0.003873,
  0.004048,   0.004048,    0.004048,    0.004048,
  0.004203,   0.004203,    0.004203,    0.004203,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004487,   0.004487,    0.004487,    0.004487,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004599,   0.004599,    0.004599,    0.004599,
  0.004642,   0.004642,    0.004642,    0.004642,
  0.0047,     0.0047,      0.0047,      0.0047,
  0.004712,   0.004712,    0.004712,    0.004712,
  0.004678,   0.004678,    0.004678,    0.004678,
  0.004661,   0.004661,    0.004661,    0.004661,
  0.004664,   0.004664,    0.004664,    0.004664,
  0.004683,   0.004683,    0.004683,    0.004683,
  0.0047,     0.0047,      0.0047,      0.0047,
  0.0047,     0.0047,      0.0047,      0.0047,
  0.0047,     0.0047,      0.0047,      0.0047,
  0.004683,   0.004683,    0.004683,    0.004683,
  0.004666,   0.004666,    0.004666,    0.004666,
  0.004666,   0.004666,    0.004666,    0.004666,
  0.004666,   0.004666,    0.004666,    0.004666,
  0.00468,    0.00468,     0.00468,     0.00468,
  0.004712,   0.004712,    0.004712,    0.004712,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004773,   0.004773,    0.004773,    0.004773,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004773,   0.004773,    0.004773,    0.004773,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004773,   0.004773,    0.004773,    0.004773,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.005045,   0.005045,    0.005045,    0.005045,
  0.005234,   0.005234,    0.005234,    0.005234,
  0.005365,   0.005365,    0.005365,    0.005365,
  0.005489,   0.005489,    0.005489,    0.005489,
  0.005671,   0.005671,    0.005671,    0.005671,
  0.005685,   0.005685,    0.005685,    0.005685,
  0.005641,   0.005641,    0.005641,    0.005641,
  0.005672,   0.005672,    0.005672,    0.005672,
  0.005643,   0.005643,    0.005643,    0.005643,
  0.005578,   0.005578,    0.005578,    0.005578,
  0.005487,   0.005487,    0.005487,    0.005487,
  0.005312,   0.005312,    0.005312,    0.005312,
  0.005096,   0.005096,    0.005096,    0.005096,
  0.004925,   0.004925,    0.004925,    0.004925,
  0.004812,   0.004812,    0.004812,    0.004812,
  0.00479,    0.00479,     0.00479,     0.00479,
  0.0048,     0.0048,      0.0048,      0.0048,
  0.004761,   0.004761,    0.004761,    0.004761,
  0.004643,   0.004643,    0.004643,    0.004643,
  0.004492,   0.004492,    0.004492,    0.004492,
  0.004436,   0.004436,    0.004436,    0.004436,
  0.004415,   0.004415,    0.004415,    0.004415,
  0.004398,   0.004398,    0.004398,    0.004398,
  0.004319,   0.004319,    0.004319,    0.004319,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.003791,   0.003791,    0.003791,    0.003791,
  0.003578,   0.003578,    0.003578,    0.003578,
  0.00346,    0.00346,     0.00346,     0.00346,
  0.003405,   0.003405,    0.003405,    0.003405,
  0.003416,   0.003416,    0.003416,    0.003416,
  0.003409,   0.003409,    0.003409,    0.003409,
  0.003386,   0.003386,    0.003386,    0.003386,
  0.003364,   0.003364,    0.003364,    0.003364,
  0.00331,    0.00331,     0.00331,     0.00331,
  0.003257,   0.003257,    0.003257,    0.003257,
  0.003249,   0.003249,    0.003249,    0.003249,
  0.003242,   0.003242,    0.003242,    0.003242,
  0.003191,   0.003191,    0.003191,    0.003191,
  0.003089,   0.003089,    0.003089,    0.003089,
  0.002969,   0.002969,    0.002969,    0.002969,
  0.002913,   0.002913,    0.002913,    0.002913,
  0.002907,   0.002907,    0.002907,    0.002907,
  0.00292,    0.00292,     0.00292,     0.00292,
  0.002954,   0.002954,    0.002954,    0.002954,
  0.002981,   0.002981,    0.002981,    0.002981,
  0.002993,   0.002993,    0.002993,    0.002993,
  0.003022,   0.003022,    0.003022,    0.003022,
  0.003052,   0.003052,    0.003052,    0.003052,
  0.003101,   0.003101,    0.003101,    0.003101,
  0.00318,    0.00318,     0.00318,     0.00318,
  0.003229,   0.003229,    0.003229,    0.003229,
  0.003265,   0.003265,    0.003265,    0.003265,
  0.003312,   0.003312,    0.003312,    0.003312,
  0.003336,   0.003336,    0.003336,    0.003336,
  0.003331,   0.003331,    0.003331,    0.003331,
  0.003344,   0.003344,    0.003344,    0.003344,
  0.003377,   0.003377,    0.003377,    0.003377,
  0.003391,   0.003391,    0.003391,    0.003391,
  0.003414,   0.003414,    0.003414,    0.003414,
  0.003401,   0.003401,    0.003401,    0.003401,
  0.003364,   0.003364,    0.003364,    0.003364,
  0.003399,   0.003399,    0.003399,    0.003399,
  0.00346,    0.00346,     0.00346,     0.00346,
  0.003473,   0.003473,    0.003473,    0.003473,
  0.003446,   0.003446,    0.003446,    0.003446,
  0.003396,   0.003396,    0.003396,    0.003396,
  0.003363,   0.003363,    0.003363,    0.003363,
  0.003377,   0.003377,    0.003377,    0.003377,
  0.003391,   0.003391,    0.003391,    0.003391,
  0.003421,   0.003421,    0.003421,    0.003421,
  0.003453,   0.003453,    0.003453,    0.003453,
  0.003485,   0.003485,    0.003485,    0.003485,
  0.003565,   0.003565,    0.003565,    0.003565,
  0.003869,   0.003869,    0.003869,    0.003869,
  0.004252,   0.004252,    0.004252,    0.004252,
  0.004538,   0.004538,    0.004538,    0.004538,
  0.004756,   0.004756,    0.004756,    0.004756,
  0.004924,   0.004924,    0.004924,    0.004924,
  0.005076,   0.005076,    0.005076,    0.005076,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005395,   0.005395,    0.005395,    0.005395,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005561,   0.005561,    0.005561,    0.005561,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005714,   0.005714,    0.005714,    0.005714,
  0.005818,   0.005818,    0.005818,    0.005818,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006178,   0.006178,    0.006178,    0.006178,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006366,   0.006366,    0.006366,    0.006366,
  0.006499,   0.006499,    0.006499,    0.006499,
  0.006636,   0.006636,    0.006636,    0.006636,
  0.006856,   0.006856,    0.006856,    0.006856,
  0.007071,   0.007071,    0.007071,    0.007071,
  0.007187,   0.007187,    0.007187,    0.007187,
  0.007296,   0.007296,    0.007296,    0.007296,
  0.007426,   0.007426,    0.007426,    0.007426,
  0.007549,   0.007549,    0.007549,    0.007549,
  0.00764,    0.00764,     0.00764,     0.00764,
  0.007588,   0.007588,    0.007588,    0.007588,
  0.007474,   0.007474,    0.007474,    0.007474,
  0.007342,   0.007342,    0.007342,    0.007342,
  0.007224,   0.007224,    0.007224,    0.007224,
  0.007287,   0.007287,    0.007287,    0.007287,
  0.007279,   0.007279,    0.007279,    0.007279,
  0.007109,   0.007109,    0.007109,    0.007109,
  0.007149,   0.007149,    0.007149,    0.007149,
  0.007298,   0.007298,    0.007298,    0.007298,
  0.007353,   0.007353,    0.007353,    0.007353,
  0.00734,    0.00734,     0.00734,     0.00734,
  0.007257,   0.007257,    0.007257,    0.007257,
  0.007148,   0.007148,    0.007148,    0.007148,
  0.007072,   0.007072,    0.007072,    0.007072,
  0.006997,   0.006997,    0.006997,    0.006997,
  0.006882,   0.006882,    0.006882,    0.006882,
  0.00679,    0.00679,     0.00679,     0.00679,
  0.006729,   0.006729,    0.006729,    0.006729,
  0.00672,    0.00672,     0.00672,     0.00672,
  0.006732,   0.006732,    0.006732,    0.006732,
  0.006761,   0.006761,    0.006761,    0.006761,
  0.006831,   0.006831,    0.006831,    0.006831,
  0.006893,   0.006893,    0.006893,    0.006893,
  0.006934,   0.006934,    0.006934,    0.006934,
  0.006934,   0.006934,    0.006934,    0.006934,
  0.006913,   0.006913,    0.006913,    0.006913,
  0.006903,   0.006903,    0.006903,    0.006903,
  0.006913,   0.006913,    0.006913,    0.006913,
  0.006944,   0.006944,    0.006944,    0.006944,
  0.006976,   0.006976,    0.006976,    0.006976,
  0.007028,   0.007028,    0.007028,    0.007028,
  0.007133,   0.007133,    0.007133,    0.007133,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007249,   0.007249,    0.007249,    0.007249,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007186,   0.007186,    0.007186,    0.007186,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.00725,    0.00725,     0.00725,     0.00725,
  0.007378,   0.007378,    0.007378,    0.007378,
  0.007544,   0.007544,    0.007544,    0.007544,
  0.007636,   0.007636,    0.007636,    0.007636,
  0.007624,   0.007624,    0.007624,    0.007624,
  0.007581,   0.007581,    0.007581,    0.007581,
  0.007516,   0.007516,    0.007516,    0.007516,
  0.007405,   0.007405,    0.007405,    0.007405,
  0.00735,    0.00735,     0.00735,     0.00735,
  0.007311,   0.007311,    0.007311,    0.007311,
  0.007233,   0.007233,    0.007233,    0.007233,
  0.007178,   0.007178,    0.007178,    0.007178,
  0.007083,   0.007083,    0.007083,    0.007083,
  0.00702,    0.00702,     0.00702,     0.00702,
  0.006989,   0.006989,    0.006989,    0.006989,
  0.006972,   0.006972,    0.006972,    0.006972,
  0.007021,   0.007021,    0.007021,    0.007021,
  0.007034,   0.007034,    0.007034,    0.007034,
  0.006977,   0.006977,    0.006977,    0.006977,
  0.006924,   0.006924,    0.006924,    0.006924,
  0.006904,   0.006904,    0.006904,    0.006904,
  0.006883,   0.006883,    0.006883,    0.006883,
  0.006904,   0.006904,    0.006904,    0.006904,
  0.006956,   0.006956,    0.006956,    0.006956,
  0.006997,   0.006997,    0.006997,    0.006997,
  0.007029,   0.007029,    0.007029,    0.007029,
  0.007039,   0.007039,    0.007039,    0.007039,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007292,   0.007292,    0.007292,    0.007292,
  0.007356,   0.007356,    0.007356,    0.007356,
  0.007335,   0.007335,    0.007335,    0.007335,
  0.007271,   0.007271,    0.007271,    0.007271,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.00725,    0.00725,     0.00725,     0.00725,
  0.007292,   0.007292,    0.007292,    0.007292,
  0.007292,   0.007292,    0.007292,    0.007292,
  0.007357,   0.007357,    0.007357,    0.007357,
  0.007554,   0.007554,    0.007554,    0.007554,
  0.007782,   0.007782,    0.007782,    0.007782,
  0.007878,   0.007878,    0.007878,    0.007878,
  0.007712,   0.007712,    0.007712,    0.007712,
  0.007445,   0.007445,    0.007445,    0.007445,
  0.007203,   0.007203,    0.007203,    0.007203,
  0.006988,   0.006988,    0.006988,    0.006988,
  0.006808,   0.006808,    0.006808,    0.006808,
  0.006724,   0.006724,    0.006724,    0.006724,
  0.006745,   0.006745,    0.006745,    0.006745,
  0.006724,   0.006724,    0.006724,    0.006724,
  0.006777,   0.006777,    0.006777,    0.006777,
  0.006861,   0.006861,    0.006861,    0.006861,
  0.006881,   0.006881,    0.006881,    0.006881,
  0.006903,   0.006903,    0.006903,    0.006903,
  0.006924,   0.006924,    0.006924,    0.006924,
  0.006935,   0.006935,    0.006935,    0.006935,
  0.006946,   0.006946,    0.006946,    0.006946,
  0.006978,   0.006978,    0.006978,    0.006978,
  0.006987,   0.006987,    0.006987,    0.006987,
  0.006976,   0.006976,    0.006976,    0.006976,
  0.007008,   0.007008,    0.007008,    0.007008,
  0.007008,   0.007008,    0.007008,    0.007008,
  0.006966,   0.006966,    0.006966,    0.006966,
  0.006944,   0.006944,    0.006944,    0.006944,
  0.006955,   0.006955,    0.006955,    0.006955,
  0.006944,   0.006944,    0.006944,    0.006944,
  0.006902,   0.006902,    0.006902,    0.006902,
  0.006913,   0.006913,    0.006913,    0.006913,
  0.006924,   0.006924,    0.006924,    0.006924,
  0.006861,   0.006861,    0.006861,    0.006861,
  0.006767,   0.006767,    0.006767,    0.006767,
  0.00663,    0.00663,     0.00663,     0.00663,
  0.006462,   0.006462,    0.006462,    0.006462,
  0.006277,   0.006277,    0.006277,    0.006277,
  0.006102,   0.006102,    0.006102,    0.006102,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006065,   0.006065,    0.006065,    0.006065,
  0.006028,   0.006028,    0.006028,    0.006028,
  0.005957,   0.005957,    0.005957,    0.005957,
  0.005957,   0.005957,    0.005957,    0.005957,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.006147,   0.006147,    0.006147,    0.006147,
  0.006183,   0.006183,    0.006183,    0.006183,
  0.006113,   0.006113,    0.006113,    0.006113,
  0.006058,   0.006058,    0.006058,    0.006058,
  0.006015,   0.006015,    0.006015,    0.006015,
  0.005983,   0.005983,    0.005983,    0.005983,
  0.005932,   0.005932,    0.005932,    0.005932,
  0.005876,   0.005876,    0.005876,    0.005876,
  0.005821,   0.005821,    0.005821,    0.005821,
  0.005722,   0.005722,    0.005722,    0.005722,
  0.005667,   0.005667,    0.005667,    0.005667,
  0.005659,   0.005659,    0.005659,    0.005659,
  0.005644,   0.005644,    0.005644,    0.005644,
  0.00566,    0.00566,     0.00566,     0.00566,
  0.005681,   0.005681,    0.005681,    0.005681,
  0.005697,   0.005697,    0.005697,    0.005697,
  0.00579,    0.00579,     0.00579,     0.00579,
  0.005907,   0.005907,    0.005907,    0.005907,
  0.00597,    0.00597,     0.00597,     0.00597,
  0.006063,   0.006063,    0.006063,    0.006063,
  0.006189,   0.006189,    0.006189,    0.006189,
  0.006253,   0.006253,    0.006253,    0.006253,
  0.006278,   0.006278,    0.006278,    0.006278,
  0.006233,   0.006233,    0.006233,    0.006233,
  0.006133,   0.006133,    0.006133,    0.006133,
  0.006084,   0.006084,    0.006084,    0.006084,
  0.00604,    0.00604,     0.00604,     0.00604,
  0.005934,   0.005934,    0.005934,    0.005934,
  0.005785,   0.005785,    0.005785,    0.005785,
  0.005734,   0.005734,    0.005734,    0.005734,
  0.005765,   0.005765,    0.005765,    0.005765,
  0.005735,   0.005735,    0.005735,    0.005735,
  0.005657,   0.005657,    0.005657,    0.005657,
  0.005614,   0.005614,    0.005614,    0.005614,
  0.005592,   0.005592,    0.005592,    0.005592,
  0.00557,    0.00557,     0.00557,     0.00557,
  0.005548,   0.005548,    0.005548,    0.005548,
  0.00552,    0.00552,     0.00552,     0.00552,
  0.005492,   0.005492,    0.005492,    0.005492,
  0.005452,   0.005452,    0.005452,    0.005452,
  0.005412,   0.005412,    0.005412,    0.005412,
  0.00536,    0.00536,     0.00536,     0.00536,
  0.005349,   0.005349,    0.005349,    0.005349,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005443,   0.005443,    0.005443,    0.005443,
  0.005579,   0.005579,    0.005579,    0.005579,
  0.005664,   0.005664,    0.005664,    0.005664,
  0.005569,   0.005569,    0.005569,    0.005569,
  0.005804,   0.005804,    0.005804,    0.005804,
  0.006286,   0.006286,    0.006286,    0.006286,
  0.006482,   0.006482,    0.006482,    0.006482,
  0.006526,   0.006526,    0.006526,    0.006526,
  0.006565,   0.006565,    0.006565,    0.006565,
  0.006561,   0.006561,    0.006561,    0.006561,
  0.006569,   0.006569,    0.006569,    0.006569,
  0.006609,   0.006609,    0.006609,    0.006609,
  0.006669,   0.006669,    0.006669,    0.006669,
  0.006709,   0.006709,    0.006709,    0.006709,
  0.006657,   0.006657,    0.006657,    0.006657,
  0.006514,   0.006514,    0.006514,    0.006514,
  0.006275,   0.006275,    0.006275,    0.006275,
  0.006139,   0.006139,    0.006139,    0.006139,
  0.006165,   0.006165,    0.006165,    0.006165,
  0.006209,   0.006209,    0.006209,    0.006209,
  0.006268,   0.006268,    0.006268,    0.006268,
  0.00624,    0.00624,     0.00624,     0.00624,
  0.00617,    0.00617,     0.00617,     0.00617,
  0.006031,   0.006031,    0.006031,    0.006031,
  0.005854,   0.005854,    0.005854,    0.005854,
  0.005764,   0.005764,    0.005764,    0.005764,
  0.005694,   0.005694,    0.005694,    0.005694,
  0.005644,   0.005644,    0.005644,    0.005644,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005499,   0.005499,    0.005499,    0.005499,
  0.005292,   0.005292,    0.005292,    0.005292,
  0.00513,    0.00513,     0.00513,     0.00513,
  0.005108,   0.005108,    0.005108,    0.005108,
  0.005116,   0.005116,    0.005116,    0.005116,
  0.005108,   0.005108,    0.005108,    0.005108,
  0.005055,   0.005055,    0.005055,    0.005055,
  0.005025,   0.005025,    0.005025,    0.005025,
  0.005112,   0.005112,    0.005112,    0.005112,
  0.005165,   0.005165,    0.005165,    0.005165,
  0.005102,   0.005102,    0.005102,    0.005102,
  0.005074,   0.005074,    0.005074,    0.005074,
  0.005081,   0.005081,    0.005081,    0.005081,
  0.005128,   0.005128,    0.005128,    0.005128,
  0.005196,   0.005196,    0.005196,    0.005196,
  0.005194,   0.005194,    0.005194,    0.005194,
  0.005162,   0.005162,    0.005162,    0.005162,
  0.005163,   0.005163,    0.005163,    0.005163,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005246,   0.005246,    0.005246,    0.005246,
  0.005271,   0.005271,    0.005271,    0.005271,
  0.005409,   0.005409,    0.005409,    0.005409,
  0.005654,   0.005654,    0.005654,    0.005654,
  0.005893,   0.005893,    0.005893,    0.005893,
  0.006006,   0.006006,    0.006006,    0.006006,
  0.005962,   0.005962,    0.005962,    0.005962,
  0.005881,   0.005881,    0.005881,    0.005881,
  0.005806,   0.005806,    0.005806,    0.005806,
  0.005706,   0.005706,    0.005706,    0.005706,
  0.00565,    0.00565,     0.00565,     0.00565,
  0.005659,   0.005659,    0.005659,    0.005659,
  0.005649,   0.005649,    0.005649,    0.005649,
  0.005595,   0.005595,    0.005595,    0.005595,
  0.00555,    0.00555,     0.00555,     0.00555,
  0.00557,    0.00557,     0.00557,     0.00557,
  0.005604,   0.005604,    0.005604,    0.005604,
  0.005622,   0.005622,    0.005622,    0.005622,
  0.005647,   0.005647,    0.005647,    0.005647,
  0.005654,   0.005654,    0.005654,    0.005654,
  0.005664,   0.005664,    0.005664,    0.005664,
  0.005699,   0.005699,    0.005699,    0.005699,
  0.005704,   0.005704,    0.005704,    0.005704,
  0.005667,   0.005667,    0.005667,    0.005667,
  0.005602,   0.005602,    0.005602,    0.005602,
  0.005516,   0.005516,    0.005516,    0.005516,
  0.005423,   0.005423,    0.005423,    0.005423,
  0.00534,    0.00534,     0.00534,     0.00534,
  0.00526,    0.00526,     0.00526,     0.00526,
  0.005113,   0.005113,    0.005113,    0.005113,
  0.00499,    0.00499,     0.00499,     0.00499,
  0.005077,   0.005077,    0.005077,    0.005077,
  0.005187,   0.005187,    0.005187,    0.005187,
  0.005081,   0.005081,    0.005081,    0.005081,
  0.004984,   0.004984,    0.004984,    0.004984,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.00533,    0.00533,     0.00533,     0.00533,
  0.005907,   0.005907,    0.005907,    0.005907,
  0.00622,    0.00622,     0.00622,     0.00622,
  0.006277,   0.006277,    0.006277,    0.006277,
  0.00629,    0.00629,     0.00629,     0.00629,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006315,   0.006315,    0.006315,    0.006315,
  0.006252,   0.006252,    0.006252,    0.006252,
  0.006164,   0.006164,    0.006164,    0.006164,
  0.006076,   0.006076,    0.006076,    0.006076,
  0.006026,   0.006026,    0.006026,    0.006026,
  0.005989,   0.005989,    0.005989,    0.005989,
  0.005929,   0.005929,    0.005929,    0.005929,
  0.005916,   0.005916,    0.005916,    0.005916,
  0.005894,   0.005894,    0.005894,    0.005894,
  0.005845,   0.005845,    0.005845,    0.005845,
  0.005769,   0.005769,    0.005769,    0.005769,
  0.005698,   0.005698,    0.005698,    0.005698,
  0.005698,   0.005698,    0.005698,    0.005698,
  0.005604,   0.005604,    0.005604,    0.005604,
  0.005478,   0.005478,    0.005478,    0.005478,
  0.005472,   0.005472,    0.005472,    0.005472,
  0.005448,   0.005448,    0.005448,    0.005448,
  0.005393,   0.005393,    0.005393,    0.005393,
  0.005366,   0.005366,    0.005366,    0.005366,
  0.005346,   0.005346,    0.005346,    0.005346,
  0.005316,   0.005316,    0.005316,    0.005316,
  0.005279,   0.005279,    0.005279,    0.005279,
  0.00526,    0.00526,     0.00526,     0.00526,
  0.005256,   0.005256,    0.005256,    0.005256,
  0.005275,   0.005275,    0.005275,    0.005275,
  0.005305,   0.005305,    0.005305,    0.005305,
  0.005326,   0.005326,    0.005326,    0.005326,
  0.005367,   0.005367,    0.005367,    0.005367,
  0.00544,    0.00544,     0.00544,     0.00544,
  0.005452,   0.005452,    0.005452,    0.005452,
  0.005439,   0.005439,    0.005439,    0.005439,
  0.005453,   0.005453,    0.005453,    0.005453,
  0.005409,   0.005409,    0.005409,    0.005409,
  0.005541,   0.005541,    0.005541,    0.005541,
  0.00579,    0.00579,     0.00579,     0.00579,
  0.00583,    0.00583,     0.00583,     0.00583,
  0.005655,   0.005655,    0.005655,    0.005655,
  0.005517,   0.005517,    0.005517,    0.005517,
  0.005529,   0.005529,    0.005529,    0.005529,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.00556,    0.00556,     0.00556,     0.00556,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005714,   0.005714,    0.005714,    0.005714,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005714,   0.005714,    0.005714,    0.005714,
  0.005714,   0.005714,    0.005714,    0.005714,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005836,   0.005836,    0.005836,    0.005836,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.005836,   0.005836,    0.005836,    0.005836,
  0.005697,   0.005697,    0.005697,    0.005697,
  0.005561,   0.005561,    0.005561,    0.005561,
  0.005444,   0.005444,    0.005444,    0.005444,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.004893,   0.004893,    0.004893,    0.004893,
  0.004773,   0.004773,    0.004773,    0.004773,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004999,   0.004999,    0.004999,    0.004999,
  0.004896,   0.004896,    0.004896,    0.004896,
  0.004714,   0.004714,    0.004714,    0.004714,
  0.004601,   0.004601,    0.004601,    0.004601,
  0.004543,   0.004543,    0.004543,    0.004543,
  0.004805,   0.004805,    0.004805,    0.004805,
  0.005045,   0.005045,    0.005045,    0.005045,
  0.005283,   0.005283,    0.005283,    0.005283,
  0.005613,   0.005613,    0.005613,    0.005613,
  0.005854,   0.005854,    0.005854,    0.005854,
  0.005996,   0.005996,    0.005996,    0.005996,
  0.006142,   0.006142,    0.006142,    0.006142,
  0.006252,   0.006252,    0.006252,    0.006252,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006142,   0.006142,    0.006142,    0.006142,
  0.005996,   0.005996,    0.005996,    0.005996,
  0.005871,   0.005871,    0.005871,    0.005871,
  0.005766,   0.005766,    0.005766,    0.005766,
  0.005697,   0.005697,    0.005697,    0.005697,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005494,   0.005494,    0.005494,    0.005494,
  0.005298,   0.005298,    0.005298,    0.005298,
  0.005107,   0.005107,    0.005107,    0.005107,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005394,   0.005394,    0.005394,    0.005394,
  0.005394,   0.005394,    0.005394,    0.005394,
  0.00533,    0.00533,     0.00533,     0.00533,
  0.00525,    0.00525,     0.00525,     0.00525,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005314,   0.005314,    0.005314,    0.005314,
  0.005316,   0.005316,    0.005316,    0.005316,
  0.005334,   0.005334,    0.005334,    0.005334,
  0.005334,   0.005334,    0.005334,    0.005334,
  0.005286,   0.005286,    0.005286,    0.005286,
  0.005206,   0.005206,    0.005206,    0.005206,
  0.005109,   0.005109,    0.005109,    0.005109,
  0.005061,   0.005061,    0.005061,    0.005061,
  0.005045,   0.005045,    0.005045,    0.005045,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.005059,   0.005059,    0.005059,    0.005059,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004877,   0.004877,    0.004877,    0.004877,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.004891,   0.004891,    0.004891,    0.004891,
  0.00483,    0.00483,     0.00483,     0.00483,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004906,   0.004906,    0.004906,    0.004906,
  0.005028,   0.005028,    0.005028,    0.005028,
  0.005145,   0.005145,    0.005145,    0.005145,
  0.005222,   0.005222,    0.005222,    0.005222,
  0.005311,   0.005311,    0.005311,    0.005311,
  0.005381,   0.005381,    0.005381,    0.005381,
  0.005398,   0.005398,    0.005398,    0.005398,
  0.005458,   0.005458,    0.005458,    0.005458,
  0.005538,   0.005538,    0.005538,    0.005538,
  0.005609,   0.005609,    0.005609,    0.005609,
  0.005663,   0.005663,    0.005663,    0.005663,
  0.005631,   0.005631,    0.005631,    0.005631,
  0.0056,     0.0056,      0.0056,      0.0056,
  0.005636,   0.005636,    0.005636,    0.005636,
  0.005636,   0.005636,    0.005636,    0.005636,
  0.005649,   0.005649,    0.005649,    0.005649,
  0.005681,   0.005681,    0.005681,    0.005681,
  0.005681,   0.005681,    0.005681,    0.005681,
  0.005694,   0.005694,    0.005694,    0.005694,
  0.005708,   0.005708,    0.005708,    0.005708,
  0.005651,   0.005651,    0.005651,    0.005651,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005522,   0.005522,    0.005522,    0.005522,
  0.005485,   0.005485,    0.005485,    0.005485,
  0.005522,   0.005522,    0.005522,    0.005522,
  0.005566,   0.005566,    0.005566,    0.005566,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005595,   0.005595,    0.005595,    0.005595,
  0.005582,   0.005582,    0.005582,    0.005582,
  0.005582,   0.005582,    0.005582,    0.005582,
  0.005555,   0.005555,    0.005555,    0.005555,
  0.005533,   0.005533,    0.005533,    0.005533,
  0.005582,   0.005582,    0.005582,    0.005582,
  0.005614,   0.005614,    0.005614,    0.005614,
  0.005659,   0.005659,    0.005659,    0.005659,
  0.005744,   0.005744,    0.005744,    0.005744,
  0.005784,   0.005784,    0.005784,    0.005784,
  0.005826,   0.005826,    0.005826,    0.005826,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.005978,   0.005978,    0.005978,    0.005978,
  0.006032,   0.006032,    0.006032,    0.006032,
  0.006086,   0.006086,    0.006086,    0.006086,
  0.006123,   0.006123,    0.006123,    0.006123,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.006197,   0.006197,    0.006197,    0.006197,
  0.006252,   0.006252,    0.006252,    0.006252,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006422,   0.006422,    0.006422,    0.006422,
  0.006461,   0.006461,    0.006461,    0.006461,
  0.006519,   0.006519,    0.006519,    0.006519,
  0.006577,   0.006577,    0.006577,    0.006577,
  0.006636,   0.006636,    0.006636,    0.006636,
  0.006715,   0.006715,    0.006715,    0.006715,
  0.006775,   0.006775,    0.006775,    0.006775,
  0.006815,   0.006815,    0.006815,    0.006815,
  0.006835,   0.006835,    0.006835,    0.006835,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006875,   0.006875,    0.006875,    0.006875,
  0.006896,   0.006896,    0.006896,    0.006896,
  0.006937,   0.006937,    0.006937,    0.006937,
  0.006978,   0.006978,    0.006978,    0.006978,
  0.006998,   0.006998,    0.006998,    0.006998,
  0.006998,   0.006998,    0.006998,    0.006998,
  0.007019,   0.007019,    0.007019,    0.007019,
  0.007039,   0.007039,    0.007039,    0.007039,
  0.007039,   0.007039,    0.007039,    0.007039,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007249,   0.007249,    0.007249,    0.007249,
  0.007249,   0.007249,    0.007249,    0.007249,
  0.007228,   0.007228,    0.007228,    0.007228,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007186,   0.007186,    0.007186,    0.007186,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007154,   0.007154,    0.007154,    0.007154,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007134,   0.007134,    0.007134,    0.007134,
  0.007134,   0.007134,    0.007134,    0.007134,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007039,   0.007039,    0.007039,    0.007039,
  0.006977,   0.006977,    0.006977,    0.006977,
  0.006915,   0.006915,    0.006915,    0.006915,
  0.006813,   0.006813,    0.006813,    0.006813,
  0.006672,   0.006672,    0.006672,    0.006672,
  0.006502,   0.006502,    0.006502,    0.006502,
  0.006354,   0.006354,    0.006354,    0.006354,
  0.006277,   0.006277,    0.006277,    0.006277,
  0.006258,   0.006258,    0.006258,    0.006258,
  0.00622,    0.00622,     0.00622,     0.00622,
  0.006158,   0.006158,    0.006158,    0.006158,
  0.006102,   0.006102,    0.006102,    0.006102,
  0.005934,   0.005934,    0.005934,    0.005934,
  0.005776,   0.005776,    0.005776,    0.005776,
  0.005693,   0.005693,    0.005693,    0.005693,
  0.005583,   0.005583,    0.005583,    0.005583,
  0.005448,   0.005448,    0.005448,    0.005448,
  0.0053,     0.0053,      0.0053,      0.0053,
  0.005187,   0.005187,    0.005187,    0.005187,
  0.005108,   0.005108,    0.005108,    0.005108,
  0.005061,   0.005061,    0.005061,    0.005061,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.004982,   0.004982,    0.004982,    0.004982,
  0.004981,   0.004981,    0.004981,    0.004981,
  0.004981,   0.004981,    0.004981,    0.004981,
  0.004933,   0.004933,    0.004933,    0.004933,
  0.004886,   0.004886,    0.004886,    0.004886,
  0.00484,    0.00484,     0.00484,     0.00484,
  0.00481,    0.00481,     0.00481,     0.00481,
  0.004811,   0.004811,    0.004811,    0.004811,
  0.004811,   0.004811,    0.004811,    0.004811,
  0.00478,    0.00478,     0.00478,     0.00478,
  0.004762,   0.004762,    0.004762,    0.004762,
  0.00476,    0.00476,     0.00476,     0.00476,
  0.004777,   0.004777,    0.004777,    0.004777,
  0.004831,   0.004831,    0.004831,    0.004831,
  0.00487,    0.00487,     0.00487,     0.00487,
  0.004927,   0.004927,    0.004927,    0.004927,
  0.004989,   0.004989,    0.004989,    0.004989,
  0.004985,   0.004985,    0.004985,    0.004985,
  0.004948,   0.004948,    0.004948,    0.004948,
  0.004916,   0.004916,    0.004916,    0.004916,
  0.004809,   0.004809,    0.004809,    0.004809,
  0.004734,   0.004734,    0.004734,    0.004734,
  0.004722,   0.004722,    0.004722,    0.004722,
  0.004819,   0.004819,    0.004819,    0.004819,
  0.004935,   0.004935,    0.004935,    0.004935,
  0.004884,   0.004884,    0.004884,    0.004884,
  0.004841,   0.004841,    0.004841,    0.004841,
  0.00488,    0.00488,     0.00488,     0.00488,
  0.004893,   0.004893,    0.004893,    0.004893,
  0.004875,   0.004875,    0.004875,    0.004875,
  0.004841,   0.004841,    0.004841,    0.004841,
  0.004823,   0.004823,    0.004823,    0.004823,
  0.004808,   0.004808,    0.004808,    0.004808,
  0.00473,    0.00473,     0.00473,     0.00473,
  0.004652,   0.004652,    0.004652,    0.004652,
  0.004576,   0.004576,    0.004576,    0.004576,
  0.004454,   0.004454,    0.004454,    0.004454,
  0.004347,   0.004347,    0.004347,    0.004347,
  0.004273,   0.004273,    0.004273,    0.004273,
  0.004218,   0.004218,    0.004218,    0.004218,
  0.004168,   0.004168,    0.004168,    0.004168,
  0.00412,    0.00412,     0.00412,     0.00412,
  0.004102,   0.004102,    0.004102,    0.004102,
  0.004053,   0.004053,    0.004053,    0.004053,
  0.004,      0.004,       0.004,       0.004,
  0.003987,   0.003987,    0.003987,    0.003987,
  0.004018,   0.004018,    0.004018,    0.004018,
  0.004032,   0.004032,    0.004032,    0.004032,
  0.004026,   0.004026,    0.004026,    0.004026,
  0.004066,   0.004066,    0.004066,    0.004066,
  0.004106,   0.004106,    0.004106,    0.004106,
  0.004106,   0.004106,    0.004106,    0.004106,
  0.004093,   0.004093,    0.004093,    0.004093,
  0.004106,   0.004106,    0.004106,    0.004106,
  0.004106,   0.004106,    0.004106,    0.004106,
  0.004079,   0.004079,    0.004079,    0.004079,
  0.004106,   0.004106,    0.004106,    0.004106,
  0.004138,   0.004138,    0.004138,    0.004138,
  0.004134,   0.004134,    0.004134,    0.004134,
  0.004161,   0.004161,    0.004161,    0.004161,
  0.004165,   0.004165,    0.004165,    0.004165,
  0.004178,   0.004178,    0.004178,    0.004178,
  0.004214,   0.004214,    0.004214,    0.004214,
  0.004204,   0.004204,    0.004204,    0.004204,
  0.004211,   0.004211,    0.004211,    0.004211,
  0.004254,   0.004254,    0.004254,    0.004254,
  0.004286,   0.004286,    0.004286,    0.004286,
  0.004336,   0.004336,    0.004336,    0.004336,
  0.004351,   0.004351,    0.004351,    0.004351,
  0.004344,   0.004344,    0.004344,    0.004344,
  0.004394,   0.004394,    0.004394,    0.004394,
  0.004433,   0.004433,    0.004433,    0.004433,
  0.004475,   0.004475,    0.004475,    0.004475,
  0.004545,   0.004545,    0.004545,    0.004545,
  0.004591,   0.004591,    0.004591,    0.004591,
  0.004584,   0.004584,    0.004584,    0.004584,
  0.004515,   0.004515,    0.004515,    0.004515,
  0.004448,   0.004448,    0.004448,    0.004448,
  0.00443,    0.00443,     0.00443,     0.00443,
  0.004447,   0.004447,    0.004447,    0.004447,
  0.004433,   0.004433,    0.004433,    0.004433,
  0.004373,   0.004373,    0.004373,    0.004373,
  0.004313,   0.004313,    0.004313,    0.004313,
  0.004269,   0.004269,    0.004269,    0.004269,
  0.004225,   0.004225,    0.004225,    0.004225,
  0.004213,   0.004213,    0.004213,    0.004213,
  0.004201,   0.004201,    0.004201,    0.004201,
  0.004161,   0.004161,    0.004161,    0.004161,
  0.004168,   0.004168,    0.004168,    0.004168,
  0.004158,   0.004158,    0.004158,    0.004158,
  0.004134,   0.004134,    0.004134,    0.004134,
  0.004134,   0.004134,    0.004134,    0.004134,
  0.004109,   0.004109,    0.004109,    0.004109,
  0.004084,   0.004084,    0.004084,    0.004084,
  0.004049,   0.004049,    0.004049,    0.004049,
  0.004015,   0.004015,    0.004015,    0.004015,
  0.003969,   0.003969,    0.003969,    0.003969,
  0.003902,   0.003902,    0.003902,    0.003902,
  0.003846,   0.003846,    0.003846,    0.003846,
  0.003799,   0.003799,    0.003799,    0.003799,
  0.003732,   0.003732,    0.003732,    0.003732,
  0.003644,   0.003644,    0.003644,    0.003644,
  0.003594,   0.003594,    0.003594,    0.003594,
  0.003563,   0.003563,    0.003563,    0.003563,
  0.003549,   0.003549,    0.003549,    0.003549,
  0.003511,   0.003511,    0.003511,    0.003511,
  0.003448,   0.003448,    0.003448,    0.003448,
  0.003412,   0.003412,    0.003412,    0.003412,
  0.003379,   0.003379,    0.003379,    0.003379,
  0.003355,   0.003355,    0.003355,    0.003355,
  0.003353,   0.003353,    0.003353,    0.003353,
  0.003334,   0.003334,    0.003334,    0.003334,
  0.003241,   0.003241,    0.003241,    0.003241,
  0.003108,   0.003108,    0.003108,    0.003108,
  0.00298,    0.00298,     0.00298,     0.00298,
  0.002902,   0.002902,    0.002902,    0.002902,
  0.002902,   0.002902,    0.002902,    0.002902,
  0.002855,   0.002855,    0.002855,    0.002855,
  0.002744,   0.002744,    0.002744,    0.002744,
  0.002649,   0.002649,    0.002649,    0.002649,
  0.002652,   0.002652,    0.002652,    0.002652,
  0.00277,    0.00277,     0.00277,     0.00277,
  0.002847,   0.002847,    0.002847,    0.002847,
  0.002849,   0.002849,    0.002849,    0.002849,
  0.002864,   0.002864,    0.002864,    0.002864,
  0.002873,   0.002873,    0.002873,    0.002873,
  0.002851,   0.002851,    0.002851,    0.002851,
  0.002803,   0.002803,    0.002803,    0.002803,
  0.002682,   0.002682,    0.002682,    0.002682,
  0.002569,   0.002569,    0.002569,    0.002569,
  0.002543,   0.002543,    0.002543,    0.002543,
  0.00258,    0.00258,     0.00258,     0.00258,
  0.002657,   0.002657,    0.002657,    0.002657,
  0.0027,     0.0027,      0.0027,      0.0027,
  0.002708,   0.002708,    0.002708,    0.002708,
  0.002724,   0.002724,    0.002724,    0.002724,
  0.002721,   0.002721,    0.002721,    0.002721,
  0.002714,   0.002714,    0.002714,    0.002714,
  0.002697,   0.002697,    0.002697,    0.002697,
  0.002677,   0.002677,    0.002677,    0.002677,
  0.002704,   0.002704,    0.002704,    0.002704,
  0.002704,   0.002704,    0.002704,    0.002704,
  0.002677,   0.002677,    0.002677,    0.002677,
  0.002693,   0.002693,    0.002693,    0.002693,
  0.002705,   0.002705,    0.002705,    0.002705,
  0.002705,   0.002705,    0.002705,    0.002705,
  0.002736,   0.002736,    0.002736,    0.002736,
  0.002748,   0.002748,    0.002748,    0.002748,
  0.002772,   0.002772,    0.002772,    0.002772,
  0.002816,   0.002816,    0.002816,    0.002816,
  0.002816,   0.002816,    0.002816,    0.002816,
  0.002977,   0.002977,    0.002977,    0.002977,
  0.003208,   0.003208,    0.003208,    0.003208,
  0.003291,   0.003291,    0.003291,    0.003291,
  0.003283,   0.003283,    0.003283,    0.003283,
  0.003229,   0.003229,    0.003229,    0.003229,
  0.00323,    0.00323,     0.00323,     0.00323,
  0.003407,   0.003407,    0.003407,    0.003407,
  0.003635,   0.003635,    0.003635,    0.003635,
  0.003771,   0.003771,    0.003771,    0.003771,
  0.003871,   0.003871,    0.003871,    0.003871,
  0.00398,    0.00398,     0.00398,     0.00398,
  0.004098,   0.004098,    0.004098,    0.004098,
  0.004182,   0.004182,    0.004182,    0.004182,
  0.004238,   0.004238,    0.004238,    0.004238,
  0.004379,   0.004379,    0.004379,    0.004379,
  0.004531,   0.004531,    0.004531,    0.004531,
  0.00462,    0.00462,     0.00462,     0.00462,
  0.004697,   0.004697,    0.004697,    0.004697,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.004935,   0.004935,    0.004935,    0.004935,
  0.004951,   0.004951,    0.004951,    0.004951,
  0.004996,   0.004996,    0.004996,    0.004996,
  0.005012,   0.005012,    0.005012,    0.005012,
  0.005027,   0.005027,    0.005027,    0.005027,
  0.005028,   0.005028,    0.005028,    0.005028,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005092,   0.005092,    0.005092,    0.005092,
  0.005108,   0.005108,    0.005108,    0.005108,
  0.00514,    0.00514,     0.00514,     0.00514,
  0.005189,   0.005189,    0.005189,    0.005189,
  0.00527,    0.00527,     0.00527,     0.00527,
  0.005269,   0.005269,    0.005269,    0.005269,
  0.005236,   0.005236,    0.005236,    0.005236,
  0.00522,    0.00522,     0.00522,     0.00522,
  0.005205,   0.005205,    0.005205,    0.005205,
  0.00529,    0.00529,     0.00529,     0.00529,
  0.005414,   0.005414,    0.005414,    0.005414,
  0.005521,   0.005521,    0.005521,    0.005521,
  0.005591,   0.005591,    0.005591,    0.005591,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005699,   0.005699,    0.005699,    0.005699,
  0.005712,   0.005712,    0.005712,    0.005712,
  0.005672,   0.005672,    0.005672,    0.005672,
  0.005619,   0.005619,    0.005619,    0.005619,
  0.005619,   0.005619,    0.005619,    0.005619,
  0.005672,   0.005672,    0.005672,    0.005672,
  0.005757,   0.005757,    0.005757,    0.005757,
  0.005874,   0.005874,    0.005874,    0.005874,
  0.005965,   0.005965,    0.005965,    0.005965,
  0.005995,   0.005995,    0.005995,    0.005995,
  0.006057,   0.006057,    0.006057,    0.006057,
  0.006139,   0.006139,    0.006139,    0.006139,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.006206,   0.006206,    0.006206,    0.006206,
  0.006258,   0.006258,    0.006258,    0.006258,
  0.006277,   0.006277,    0.006277,    0.006277,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006332,   0.006332,    0.006332,    0.006332,
  0.006325,   0.006325,    0.006325,    0.006325,
  0.006349,   0.006349,    0.006349,    0.006349,
  0.006405,   0.006405,    0.006405,    0.006405,
  0.006417,   0.006417,    0.006417,    0.006417,
  0.00641,    0.00641,     0.00641,     0.00641,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006327,   0.006327,    0.006327,    0.006327,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006234,   0.006234,    0.006234,    0.006234,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.006141,   0.006141,    0.006141,    0.006141,
  0.006123,   0.006123,    0.006123,    0.006123,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.005978,   0.005978,    0.005978,    0.005978,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.005996,   0.005996,    0.005996,    0.005996,
  0.005929,   0.005929,    0.005929,    0.005929,
  0.005879,   0.005879,    0.005879,    0.005879,
  0.005946,   0.005946,    0.005946,    0.005946,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.005889,   0.005889,    0.005889,    0.005889,
  0.005798,   0.005798,    0.005798,    0.005798,
  0.005753,   0.005753,    0.005753,    0.005753,
  0.005741,   0.005741,    0.005741,    0.005741,
  0.005717,   0.005717,    0.005717,    0.005717,
  0.005697,   0.005697,    0.005697,    0.005697,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005784,   0.005784,    0.005784,    0.005784,
  0.005848,   0.005848,    0.005848,    0.005848,
  0.005767,   0.005767,    0.005767,    0.005767,
  0.005669,   0.005669,    0.005669,    0.005669,
  0.005642,   0.005642,    0.005642,    0.005642,
  0.005674,   0.005674,    0.005674,    0.005674,
  0.005674,   0.005674,    0.005674,    0.005674,
  0.005724,   0.005724,    0.005724,    0.005724,
  0.005769,   0.005769,    0.005769,    0.005769,
  0.00579,    0.00579,     0.00579,     0.00579,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005652,   0.005652,    0.005652,    0.005652,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005396,   0.005396,    0.005396,    0.005396,
  0.005366,   0.005366,    0.005366,    0.005366,
  0.005353,   0.005353,    0.005353,    0.005353,
  0.005371,   0.005371,    0.005371,    0.005371,
  0.005388,   0.005388,    0.005388,    0.005388,
  0.005388,   0.005388,    0.005388,    0.005388,
  0.005388,   0.005388,    0.005388,    0.005388,
  0.005357,   0.005357,    0.005357,    0.005357,
  0.005262,   0.005262,    0.005262,    0.005262,
  0.005182,   0.005182,    0.005182,    0.005182,
  0.005149,   0.005149,    0.005149,    0.005149,
  0.005084,   0.005084,    0.005084,    0.005084,
  0.005034,   0.005034,    0.005034,    0.005034,
  0.005,      0.005,       0.005,       0.005,
  0.004951,   0.004951,    0.004951,    0.004951,
  0.00495,    0.00495,     0.00495,     0.00495,
  0.004997,   0.004997,    0.004997,    0.004997,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.00509,    0.00509,     0.00509,     0.00509,
  0.005059,   0.005059,    0.005059,    0.005059,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004715,   0.004715,    0.004715,    0.004715,
  0.004543,   0.004543,    0.004543,    0.004543,
  0.004377,   0.004377,    0.004377,    0.004377,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004308,   0.004308,    0.004308,    0.004308,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004176,   0.004176,    0.004176,    0.004176,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004171,   0.004171,    0.004171,    0.004171,
  0.004187,   0.004187,    0.004187,    0.004187,
  0.004233,   0.004233,    0.004233,    0.004233,
  0.004238,   0.004238,    0.004238,    0.004238,
  0.00422,    0.00422,     0.00422,     0.00422,
  0.004203,   0.004203,    0.004203,    0.004203,
  0.004199,   0.004199,    0.004199,    0.004199,
  0.004196,   0.004196,    0.004196,    0.004196,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.004182,   0.004182,    0.004182,    0.004182,
  0.004185,   0.004185,    0.004185,    0.004185,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.004197,   0.004197,    0.004197,    0.004197,
  0.004174,   0.004174,    0.004174,    0.004174,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004161,   0.004161,    0.004161,    0.004161,
  0.004187,   0.004187,    0.004187,    0.004187,
  0.004169,   0.004169,    0.004169,    0.004169,
  0.004161,   0.004161,    0.004161,    0.004161,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.004179,   0.004179,    0.004179,    0.004179,
  0.004139,   0.004139,    0.004139,    0.004139,
  0.004113,   0.004113,    0.004113,    0.004113,
  0.004113,   0.004113,    0.004113,    0.004113,
  0.004095,   0.004095,    0.004095,    0.004095,
  0.004076,   0.004076,    0.004076,    0.004076,
  0.004063,   0.004063,    0.004063,    0.004063,
  0.004037,   0.004037,    0.004037,    0.004037,
  0.004029,   0.004029,    0.004029,    0.004029,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.003997,   0.003997,    0.003997,    0.003997,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.003921,   0.003921,    0.003921,    0.003921,
  0.003927,   0.003927,    0.003927,    0.003927,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003922,   0.003922,    0.003922,    0.003922,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003897,   0.003897,    0.003897,    0.003897,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003927,   0.003927,    0.003927,    0.003927,
  0.003921,   0.003921,    0.003921,    0.003921,
  0.003933,   0.003933,    0.003933,    0.003933,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.004055,   0.004055,    0.004055,    0.004055,
  0.00405,    0.00405,     0.00405,     0.00405,
  0.00405,    0.00405,     0.00405,     0.00405,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004118,   0.004118,    0.004118,    0.004118,
  0.004139,   0.004139,    0.004139,    0.004139,
  0.004191,   0.004191,    0.004191,    0.004191,
  0.004234,   0.004234,    0.004234,    0.004234,
  0.004261,   0.004261,    0.004261,    0.004261,
  0.004321,   0.004321,    0.004321,    0.004321,
  0.004398,   0.004398,    0.004398,    0.004398,
  0.00443,    0.00443,     0.00443,     0.00443,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004446,   0.004446,    0.004446,    0.004446,
  0.004461,   0.004461,    0.004461,    0.004461,
  0.004476,   0.004476,    0.004476,    0.004476,
  0.004493,   0.004493,    0.004493,    0.004493,
  0.004465,   0.004465,    0.004465,    0.004465,
  0.004423,   0.004423,    0.004423,    0.004423,
  0.004412,   0.004412,    0.004412,    0.004412,
  0.004397,   0.004397,    0.004397,    0.004397,
  0.004368,   0.004368,    0.004368,    0.004368,
  0.004341,   0.004341,    0.004341,    0.004341,
  0.00433,    0.00433,     0.00433,     0.00433,
  0.004344,   0.004344,    0.004344,    0.004344,
  0.004385,   0.004385,    0.004385,    0.004385,
  0.004402,   0.004402,    0.004402,    0.004402,
  0.004373,   0.004373,    0.004373,    0.004373,
  0.004385,   0.004385,    0.004385,    0.004385,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.00426,    0.00426,     0.00426,     0.00426,
  0.004214,   0.004214,    0.004214,    0.004214,
  0.004219,   0.004219,    0.004219,    0.004219,
  0.004192,   0.004192,    0.004192,    0.004192,
  0.004126,   0.004126,    0.004126,    0.004126,
  0.004061,   0.004061,    0.004061,    0.004061,
  0.004028,   0.004028,    0.004028,    0.004028,
  0.004022,   0.004022,    0.004022,    0.004022,
  0.004028,   0.004028,    0.004028,    0.004028,
  0.004061,   0.004061,    0.004061,    0.004061,
  0.004074,   0.004074,    0.004074,    0.004074,
  0.004048,   0.004048,    0.004048,    0.004048,
  0.00401,    0.00401,     0.00401,     0.00401,
  0.00399,    0.00399,     0.00399,     0.00399,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.003977,   0.003977,    0.003977,    0.003977,
  0.003965,   0.003965,    0.003965,    0.003965,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.003977,   0.003977,    0.003977,    0.003977,
  0.004023,   0.004023,    0.004023,    0.004023,
  0.004108,   0.004108,    0.004108,    0.004108,
  0.004165,   0.004165,    0.004165,    0.004165,
  0.004239,   0.004239,    0.004239,    0.004239,
  0.004316,   0.004316,    0.004316,    0.004316,
  0.004397,   0.004397,    0.004397,    0.004397,
  0.004468,   0.004468,    0.004468,    0.004468,
  0.004526,   0.004526,    0.004526,    0.004526,
  0.004587,   0.004587,    0.004587,    0.004587,
  0.004618,   0.004618,    0.004618,    0.004618,
  0.004619,   0.004619,    0.004619,    0.004619,
  0.004651,   0.004651,    0.004651,    0.004651,
  0.004651,   0.004651,    0.004651,    0.004651,
  0.00462,    0.00462,     0.00462,     0.00462,
  0.00462,    0.00462,     0.00462,     0.00462,
  0.004604,   0.004604,    0.004604,    0.004604,
  0.004603,   0.004603,    0.004603,    0.004603,
  0.004603,   0.004603,    0.004603,    0.004603,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004539,   0.004539,    0.004539,    0.004539,
  0.004539,   0.004539,    0.004539,    0.004539,
  0.004539,   0.004539,    0.004539,    0.004539,
  0.004524,   0.004524,    0.004524,    0.004524,
  0.004477,   0.004477,    0.004477,    0.004477,
  0.00443,    0.00443,     0.00443,     0.00443,
  0.004432,   0.004432,    0.004432,    0.004432,
  0.004418,   0.004418,    0.004418,    0.004418,
  0.004388,   0.004388,    0.004388,    0.004388,
  0.004358,   0.004358,    0.004358,    0.004358,
  0.004343,   0.004343,    0.004343,    0.004343,
  0.004343,   0.004343,    0.004343,    0.004343,
  0.004359,   0.004359,    0.004359,    0.004359,
  0.004391,   0.004391,    0.004391,    0.004391,
  0.004421,   0.004421,    0.004421,    0.004421,
  0.004436,   0.004436,    0.004436,    0.004436,
  0.004436,   0.004436,    0.004436,    0.004436,
  0.004421,   0.004421,    0.004421,    0.004421,
  0.004406,   0.004406,    0.004406,    0.004406,
  0.004406,   0.004406,    0.004406,    0.004406,
  0.004454,   0.004454,    0.004454,    0.004454,
  0.004456,   0.004456,    0.004456,    0.004456,
  0.004424,   0.004424,    0.004424,    0.004424,
  0.004439,   0.004439,    0.004439,    0.004439,
  0.004422,   0.004422,    0.004422,    0.004422,
  0.004421,   0.004421,    0.004421,    0.004421,
  0.004436,   0.004436,    0.004436,    0.004436,
  0.004469,   0.004469,    0.004469,    0.004469,
  0.004519,   0.004519,    0.004519,    0.004519,
  0.004517,   0.004517,    0.004517,    0.004517,
  0.004481,   0.004481,    0.004481,    0.004481,
  0.004494,   0.004494,    0.004494,    0.004494,
  0.004493,   0.004493,    0.004493,    0.004493,
  0.004492,   0.004492,    0.004492,    0.004492,
  0.004508,   0.004508,    0.004508,    0.004508,
  0.004523,   0.004523,    0.004523,    0.004523,
  0.004666,   0.004666,    0.004666,    0.004666,
  0.004841,   0.004841,    0.004841,    0.004841,
  0.004921,   0.004921,    0.004921,    0.004921,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004832,   0.004832,    0.004832,    0.004832,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004862,   0.004862,    0.004862,    0.004862,
  0.004877,   0.004877,    0.004877,    0.004877,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004907,   0.004907,    0.004907,    0.004907,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004967,   0.004967,    0.004967,    0.004967,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.005494,   0.005494,    0.005494,    0.005494,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005682,   0.005682,    0.005682,    0.005682,
  0.005651,   0.005651,    0.005651,    0.005651,
  0.005665,   0.005665,    0.005665,    0.005665,
  0.005645,   0.005645,    0.005645,    0.005645,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.00568,    0.00568,     0.00568,     0.00568,
  0.005748,   0.005748,    0.005748,    0.005748,
  0.005801,   0.005801,    0.005801,    0.005801,
  0.005836,   0.005836,    0.005836,    0.005836,
  0.005907,   0.005907,    0.005907,    0.005907,
  0.005978,   0.005978,    0.005978,    0.005978,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.006252,   0.006252,    0.006252,    0.006252,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006234,   0.006234,    0.006234,    0.006234,
  0.006234,   0.006234,    0.006234,    0.006234,
  0.006252,   0.006252,    0.006252,    0.006252,
  0.006252,   0.006252,    0.006252,    0.006252,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006327,   0.006327,    0.006327,    0.006327,
  0.006327,   0.006327,    0.006327,    0.006327,
  0.006327,   0.006327,    0.006327,    0.006327,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006422,   0.006422,    0.006422,    0.006422,
  0.006461,   0.006461,    0.006461,    0.006461,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.006461,   0.006461,    0.006461,    0.006461,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.006441,   0.006441,    0.006441,    0.006441,
  0.006461,   0.006461,    0.006461,    0.006461,
  0.006499,   0.006499,    0.006499,    0.006499,
  0.006538,   0.006538,    0.006538,    0.006538,
  0.006596,   0.006596,    0.006596,    0.006596,
  0.006695,   0.006695,    0.006695,    0.006695,
  0.006763,   0.006763,    0.006763,    0.006763,
  0.006792,   0.006792,    0.006792,    0.006792,
  0.006863,   0.006863,    0.006863,    0.006863,
  0.006882,   0.006882,    0.006882,    0.006882,
  0.006861,   0.006861,    0.006861,    0.006861,
  0.006871,   0.006871,    0.006871,    0.006871,
  0.006808,   0.006808,    0.006808,    0.006808,
  0.006745,   0.006745,    0.006745,    0.006745,
  0.006682,   0.006682,    0.006682,    0.006682,
  0.006598,   0.006598,    0.006598,    0.006598,
  0.006556,   0.006556,    0.006556,    0.006556,
  0.006567,   0.006567,    0.006567,    0.006567,
  0.006598,   0.006598,    0.006598,    0.006598,
  0.006598,   0.006598,    0.006598,    0.006598,
  0.006578,   0.006578,    0.006578,    0.006578,
  0.006557,   0.006557,    0.006557,    0.006557,
  0.006516,   0.006516,    0.006516,    0.006516,
  0.006475,   0.006475,    0.006475,    0.006475,
  0.006455,   0.006455,    0.006455,    0.006455,
  0.006457,   0.006457,    0.006457,    0.006457,
  0.00644,    0.00644,     0.00644,     0.00644,
  0.0064,     0.0064,      0.0064,      0.0064,
  0.006348,   0.006348,    0.006348,    0.006348,
  0.006277,   0.006277,    0.006277,    0.006277,
  0.006231,   0.006231,    0.006231,    0.006231,
  0.006216,   0.006216,    0.006216,    0.006216,
  0.00619,    0.00619,     0.00619,     0.00619,
  0.006164,   0.006164,    0.006164,    0.006164,
  0.006183,   0.006183,    0.006183,    0.006183,
  0.00617,    0.00617,     0.00617,     0.00617,
  0.00617,    0.00617,     0.00617,     0.00617,
  0.006189,   0.006189,    0.006189,    0.006189,
  0.006158,   0.006158,    0.006158,    0.006158,
  0.006126,   0.006126,    0.006126,    0.006126,
  0.006107,   0.006107,    0.006107,    0.006107,
  0.006069,   0.006069,    0.006069,    0.006069,
  0.006012,   0.006012,    0.006012,    0.006012,
  0.006006,   0.006006,    0.006006,    0.006006,
  0.006038,   0.006038,    0.006038,    0.006038,
  0.006006,   0.006006,    0.006006,    0.006006,
  0.005962,   0.005962,    0.005962,    0.005962,
  0.005949,   0.005949,    0.005949,    0.005949,
  0.005931,   0.005931,    0.005931,    0.005931,
  0.005943,   0.005943,    0.005943,    0.005943,
  0.005962,   0.005962,    0.005962,    0.005962,
  0.005981,   0.005981,    0.005981,    0.005981,
  0.006025,   0.006025,    0.006025,    0.006025,
  0.006057,   0.006057,    0.006057,    0.006057,
  0.006107,   0.006107,    0.006107,    0.006107,
  0.006151,   0.006151,    0.006151,    0.006151,
  0.006151,   0.006151,    0.006151,    0.006151,
  0.006138,   0.006138,    0.006138,    0.006138,
  0.006157,   0.006157,    0.006157,    0.006157,
  0.006157,   0.006157,    0.006157,    0.006157,
  0.00617,    0.00617,     0.00617,     0.00617,
  0.006214,   0.006214,    0.006214,    0.006214,
  0.006239,   0.006239,    0.006239,    0.006239,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.00629,    0.00629,     0.00629,     0.00629,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006252,   0.006252,    0.006252,    0.006252,
  0.006234,   0.006234,    0.006234,    0.006234,
  0.006215,   0.006215,    0.006215,    0.006215,
  0.006165,   0.006165,    0.006165,    0.006165,
  0.006097,   0.006097,    0.006097,    0.006097,
  0.006037,   0.006037,    0.006037,    0.006037,
  0.005838,   0.005838,    0.005838,    0.005838,
  0.005545,   0.005545,    0.005545,    0.005545,
  0.005314,   0.005314,    0.005314,    0.005314,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.004965,   0.004965,    0.004965,    0.004965,
  0.004814,   0.004814,    0.004814,    0.004814,
  0.004652,   0.004652,    0.004652,    0.004652,
  0.00454,    0.00454,     0.00454,     0.00454,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.00421,    0.00421,     0.00421,     0.00421,
  0.004165,   0.004165,    0.004165,    0.004165,
  0.004139,   0.004139,    0.004139,    0.004139,
  0.004093,   0.004093,    0.004093,    0.004093,
  0.004111,   0.004111,    0.004111,    0.004111,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004067,   0.004067,    0.004067,    0.004067,
  0.003978,   0.003978,    0.003978,    0.003978,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.004068,   0.004068,    0.004068,    0.004068,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004384,   0.004384,    0.004384,    0.004384,
  0.004516,   0.004516,    0.004516,    0.004516,
  0.004527,   0.004527,    0.004527,    0.004527,
  0.004442,   0.004442,    0.004442,    0.004442,
  0.004342,   0.004342,    0.004342,    0.004342,
  0.004323,   0.004323,    0.004323,    0.004323,
  0.004383,   0.004383,    0.004383,    0.004383,
  0.004391,   0.004391,    0.004391,    0.004391,
  0.004384,   0.004384,    0.004384,    0.004384,
  0.004452,   0.004452,    0.004452,    0.004452,
  0.004496,   0.004496,    0.004496,    0.004496,
  0.004524,   0.004524,    0.004524,    0.004524,
  0.004556,   0.004556,    0.004556,    0.004556,
  0.004546,   0.004546,    0.004546,    0.004546,
  0.00448,    0.00448,     0.00448,     0.00448,
  0.004399,   0.004399,    0.004399,    0.004399,
  0.004323,   0.004323,    0.004323,    0.004323,
  0.004286,   0.004286,    0.004286,    0.004286,
  0.004264,   0.004264,    0.004264,    0.004264,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004336,   0.004336,    0.004336,    0.004336,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004098,   0.004098,    0.004098,    0.004098,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003922,   0.003922,    0.003922,    0.003922,
  0.003922,   0.003922,    0.003922,    0.003922,
  0.003922,   0.003922,    0.003922,    0.003922,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003909,   0.003909,    0.003909,    0.003909,
  0.003946,   0.003946,    0.003946,    0.003946,
  0.003972,   0.003972,    0.003972,    0.003972,
  0.003916,   0.003916,    0.003916,    0.003916,
  0.003837,   0.003837,    0.003837,    0.003837,
  0.003783,   0.003783,    0.003783,    0.003783,
  0.003746,   0.003746,    0.003746,    0.003746,
  0.003737,   0.003737,    0.003737,    0.003737,
  0.003701,   0.003701,    0.003701,    0.003701,
  0.003656,   0.003656,    0.003656,    0.003656,
  0.003642,   0.003642,    0.003642,    0.003642,
  0.00366,    0.00366,     0.00366,     0.00366,
  0.003683,   0.003683,    0.003683,    0.003683,
  0.003675,   0.003675,    0.003675,    0.003675,
  0.003693,   0.003693,    0.003693,    0.003693,
  0.003724,   0.003724,    0.003724,    0.003724,
  0.003743,   0.003743,    0.003743,    0.003743,
  0.00378,    0.00378,     0.00378,     0.00378,
  0.003816,   0.003816,    0.003816,    0.003816,
  0.003809,   0.003809,    0.003809,    0.003809,
  0.003789,   0.003789,    0.003789,    0.003789,
  0.003814,   0.003814,    0.003814,    0.003814,
  0.00382,    0.00382,     0.00382,     0.00382,
  0.003821,   0.003821,    0.003821,    0.003821,
  0.003834,   0.003834,    0.003834,    0.003834,
  0.003809,   0.003809,    0.003809,    0.003809,
  0.003797,   0.003797,    0.003797,    0.003797,
  0.003834,   0.003834,    0.003834,    0.003834,
  0.003871,   0.003871,    0.003871,    0.003871,
  0.003852,   0.003852,    0.003852,    0.003852,
  0.00382,    0.00382,     0.00382,     0.00382,
  0.003839,   0.003839,    0.003839,    0.003839,
  0.003802,   0.003802,    0.003802,    0.003802,
  0.003771,   0.003771,    0.003771,    0.003771,
  0.003789,   0.003789,    0.003789,    0.003789,
  0.003782,   0.003782,    0.003782,    0.003782,
  0.003757,   0.003757,    0.003757,    0.003757,
  0.003739,   0.003739,    0.003739,    0.003739,
  0.003722,   0.003722,    0.003722,    0.003722,
  0.003693,   0.003693,    0.003693,    0.003693,
  0.003665,   0.003665,    0.003665,    0.003665,
  0.003626,   0.003626,    0.003626,    0.003626,
  0.003566,   0.003566,    0.003566,    0.003566,
  0.003498,   0.003498,    0.003498,    0.003498,
  0.003465,   0.003465,    0.003465,    0.003465,
  0.003465,   0.003465,    0.003465,    0.003465,
  0.003476,   0.003476,    0.003476,    0.003476,
  0.003487,   0.003487,    0.003487,    0.003487,
  0.003498,   0.003498,    0.003498,    0.003498,
  0.003543,   0.003543,    0.003543,    0.003543,
  0.003658,   0.003658,    0.003658,    0.003658,
  0.003825,   0.003825,    0.003825,    0.003825,
  0.004049,   0.004049,    0.004049,    0.004049,
  0.00424,    0.00424,     0.00424,     0.00424,
  0.004259,   0.004259,    0.004259,    0.004259,
  0.004196,   0.004196,    0.004196,    0.004196,
  0.004165,   0.004165,    0.004165,    0.004165,
  0.004137,   0.004137,    0.004137,    0.004137,
  0.003971,   0.003971,    0.003971,    0.003971,
  0.003792,   0.003792,    0.003792,    0.003792,
  0.003829,   0.003829,    0.003829,    0.003829,
  0.003755,   0.003755,    0.003755,    0.003755,
  0.0035,     0.0035,      0.0035,      0.0035,
  0.003386,   0.003386,    0.003386,    0.003386,
  0.003395,   0.003395,    0.003395,    0.003395,
  0.003589,   0.003589,    0.003589,    0.003589,
  0.003917,   0.003917,    0.003917,    0.003917,
  0.00407,    0.00407,     0.00407,     0.00407,
  0.004052,   0.004052,    0.004052,    0.004052,
  0.004025,   0.004025,    0.004025,    0.004025,
  0.004061,   0.004061,    0.004061,    0.004061,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004156,   0.004156,    0.004156,    0.004156,
  0.004187,   0.004187,    0.004187,    0.004187,
  0.004219,   0.004219,    0.004219,    0.004219,
  0.00425,    0.00425,     0.00425,     0.00425,
  0.004264,   0.004264,    0.004264,    0.004264,
  0.004219,   0.004219,    0.004219,    0.004219,
  0.004158,   0.004158,    0.004158,    0.004158,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.003947,   0.003947,    0.003947,    0.003947,
  0.003872,   0.003872,    0.003872,    0.003872,
  0.00386,    0.00386,     0.00386,     0.00386,
  0.003897,   0.003897,    0.003897,    0.003897,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.003959,   0.003959,    0.003959,    0.003959,
  0.003996,   0.003996,    0.003996,    0.003996,
  0.00406,    0.00406,     0.00406,     0.00406,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.00421,    0.00421,     0.00421,     0.00421,
  0.004184,   0.004184,    0.004184,    0.004184,
  0.004229,   0.004229,    0.004229,    0.004229,
  0.004264,   0.004264,    0.004264,    0.004264,
  0.00425,    0.00425,     0.00425,     0.00425,
  0.00421,    0.00421,     0.00421,     0.00421,
  0.004161,   0.004161,    0.004161,    0.004161,
  0.00413,    0.00413,     0.00413,     0.00413,
  0.004116,   0.004116,    0.004116,    0.004116,
  0.004089,   0.004089,    0.004089,    0.004089,
  0.004075,   0.004075,    0.004075,    0.004075,
  0.004075,   0.004075,    0.004075,    0.004075,
  0.004061,   0.004061,    0.004061,    0.004061,
  0.003989,   0.003989,    0.003989,    0.003989,
  0.00393,    0.00393,     0.00393,     0.00393,
  0.003935,   0.003935,    0.003935,    0.003935,
  0.003919,   0.003919,    0.003919,    0.003919,
  0.003878,   0.003878,    0.003878,    0.003878,
  0.003846,   0.003846,    0.003846,    0.003846,
  0.003769,   0.003769,    0.003769,    0.003769,
  0.003669,   0.003669,    0.003669,    0.003669,
  0.003623,   0.003623,    0.003623,    0.003623,
  0.003623,   0.003623,    0.003623,    0.003623,
  0.003544,   0.003544,    0.003544,    0.003544,
  0.003442,   0.003442,    0.003442,    0.003442,
  0.003442,   0.003442,    0.003442,    0.003442,
  0.003421,   0.003421,    0.003421,    0.003421,
  0.003366,   0.003366,    0.003366,    0.003366,
  0.003281,   0.003281,    0.003281,    0.003281,
  0.003146,   0.003146,    0.003146,    0.003146,
  0.003188,   0.003188,    0.003188,    0.003188,
  0.003188,   0.003188,    0.003188,    0.003188,
  0.003007,   0.003007,    0.003007,    0.003007,
  0.002919,   0.002919,    0.002919,    0.002919,
  0.002939,   0.002939,    0.002939,    0.002939,
  0.002977,   0.002977,    0.002977,    0.002977,
  0.003016,   0.003016,    0.003016,    0.003016,
  0.003075,   0.003075,    0.003075,    0.003075,
  0.003115,   0.003115,    0.003115,    0.003115,
  0.003115,   0.003115,    0.003115,    0.003115,
  0.003136,   0.003136,    0.003136,    0.003136,
  0.003229,   0.003229,    0.003229,    0.003229,
  0.003334,   0.003334,    0.003334,    0.003334,
  0.003421,   0.003421,    0.003421,    0.003421,
  0.003476,   0.003476,    0.003476,    0.003476,
  0.003509,   0.003509,    0.003509,    0.003509,
  0.003509,   0.003509,    0.003509,    0.003509,
  0.003498,   0.003498,    0.003498,    0.003498,
  0.003532,   0.003532,    0.003532,    0.003532,
  0.0036,     0.0036,      0.0036,      0.0036,
  0.003693,   0.003693,    0.003693,    0.003693,
  0.0038,     0.0038,      0.0038,      0.0038,
  0.003885,   0.003885,    0.003885,    0.003885,
  0.003997,   0.003997,    0.003997,    0.003997,
  0.004093,   0.004093,    0.004093,    0.004093,
  0.004121,   0.004121,    0.004121,    0.004121,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004226,   0.004226,    0.004226,    0.004226,
  0.004344,   0.004344,    0.004344,    0.004344,
  0.00437,    0.00437,     0.00437,     0.00437,
  0.004399,   0.004399,    0.004399,    0.004399,
  0.004433,   0.004433,    0.004433,    0.004433,
  0.00447,    0.00447,     0.00447,     0.00447,
  0.004487,   0.004487,    0.004487,    0.004487,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004402,   0.004402,    0.004402,    0.004402,
  0.004347,   0.004347,    0.004347,    0.004347,
  0.004319,   0.004319,    0.004319,    0.004319,
  0.004278,   0.004278,    0.004278,    0.004278,
  0.004175,   0.004175,    0.004175,    0.004175,
  0.004118,   0.004118,    0.004118,    0.004118,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004105,   0.004105,    0.004105,    0.004105,
  0.00408,    0.00408,     0.00408,     0.00408,
  0.004047,   0.004047,    0.004047,    0.004047,
  0.004009,   0.004009,    0.004009,    0.004009,
  0.003965,   0.003965,    0.003965,    0.003965,
  0.003933,   0.003933,    0.003933,    0.003933,
  0.003889,   0.003889,    0.003889,    0.003889,
  0.003795,   0.003795,    0.003795,    0.003795,
  0.003738,   0.003738,    0.003738,    0.003738,
  0.0037,     0.0037,      0.0037,      0.0037,
  0.00365,    0.00365,     0.00365,     0.00365,
  0.003626,   0.003626,    0.003626,    0.003626,
  0.003588,   0.003588,    0.003588,    0.003588,
  0.003563,   0.003563,    0.003563,    0.003563,
  0.00355,    0.00355,     0.00355,     0.00355,
  0.0035,     0.0035,      0.0035,      0.0035,
  0.003462,   0.003462,    0.003462,    0.003462,
  0.003451,   0.003451,    0.003451,    0.003451,
  0.003478,   0.003478,    0.003478,    0.003478,
  0.003491,   0.003491,    0.003491,    0.003491,
  0.003423,   0.003423,    0.003423,    0.003423,
  0.003355,   0.003355,    0.003355,    0.003355,
  0.003305,   0.003305,    0.003305,    0.003305,
  0.003256,   0.003256,    0.003256,    0.003256,
  0.003269,   0.003269,    0.003269,    0.003269,
  0.003282,   0.003282,    0.003282,    0.003282,
  0.003292,   0.003292,    0.003292,    0.003292,
  0.003386,   0.003386,    0.003386,    0.003386,
  0.003571,   0.003571,    0.003571,    0.003571,
  0.003697,   0.003697,    0.003697,    0.003697,
  0.003755,   0.003755,    0.003755,    0.003755,
  0.003872,   0.003872,    0.003872,    0.003872,
  0.003972,   0.003972,    0.003972,    0.003972,
  0.004035,   0.004035,    0.004035,    0.004035,
  0.004124,   0.004124,    0.004124,    0.004124,
  0.004227,   0.004227,    0.004227,    0.004227,
  0.004327,   0.004327,    0.004327,    0.004327,
  0.00442,    0.00442,     0.00442,     0.00442,
  0.004473,   0.004473,    0.004473,    0.004473,
  0.004548,   0.004548,    0.004548,    0.004548,
  0.004608,   0.004608,    0.004608,    0.004608,
  0.004654,   0.004654,    0.004654,    0.004654,
  0.0047,     0.0047,      0.0047,      0.0047,
  0.004744,   0.004744,    0.004744,    0.004744,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005202,   0.005202,    0.005202,    0.005202,
  0.005218,   0.005218,    0.005218,    0.005218,
  0.005218,   0.005218,    0.005218,    0.005218,
  0.005234,   0.005234,    0.005234,    0.005234,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005218,   0.005218,    0.005218,    0.005218,
  0.005187,   0.005187,    0.005187,    0.005187,
  0.005203,   0.005203,    0.005203,    0.005203,
  0.005156,   0.005156,    0.005156,    0.005156,
  0.005012,   0.005012,    0.005012,    0.005012,
  0.004827,   0.004827,    0.004827,    0.004827,
  0.004633,   0.004633,    0.004633,    0.004633,
  0.004516,   0.004516,    0.004516,    0.004516,
  0.004502,   0.004502,    0.004502,    0.004502,
  0.004499,   0.004499,    0.004499,    0.004499,
  0.004482,   0.004482,    0.004482,    0.004482,
  0.004482,   0.004482,    0.004482,    0.004482,
  0.004482,   0.004482,    0.004482,    0.004482,
  0.004482,   0.004482,    0.004482,    0.004482,
  0.004436,   0.004436,    0.004436,    0.004436,
  0.00433,    0.00433,     0.00433,     0.00433,
  0.004231,   0.004231,    0.004231,    0.004231,
  0.004156,   0.004156,    0.004156,    0.004156,
  0.004116,   0.004116,    0.004116,    0.004116,
  0.004131,   0.004131,    0.004131,    0.004131,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.004427,   0.004427,    0.004427,    0.004427,
  0.004451,   0.004451,    0.004451,    0.004451,
  0.00449,    0.00449,     0.00449,     0.00449,
  0.004487,   0.004487,    0.004487,    0.004487,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004388,   0.004388,    0.004388,    0.004388,
  0.004329,   0.004329,    0.004329,    0.004329,
  0.004256,   0.004256,    0.004256,    0.004256,
  0.004201,   0.004201,    0.004201,    0.004201,
  0.004156,   0.004156,    0.004156,    0.004156,
  0.004057,   0.004057,    0.004057,    0.004057,
  0.003972,   0.003972,    0.003972,    0.003972,
  0.003902,   0.003902,    0.003902,    0.003902,
  0.003821,   0.003821,    0.003821,    0.003821,
  0.003788,   0.003788,    0.003788,    0.003788,
  0.003773,   0.003773,    0.003773,    0.003773,
  0.003715,   0.003715,    0.003715,    0.003715,
  0.003602,   0.003602,    0.003602,    0.003602,
  0.003481,   0.003481,    0.003481,    0.003481,
  0.003396,   0.003396,    0.003396,    0.003396,
  0.003319,   0.003319,    0.003319,    0.003319,
  0.003211,   0.003211,    0.003211,    0.003211,
  0.00313,    0.00313,     0.00313,     0.00313,
  0.003041,   0.003041,    0.003041,    0.003041,
  0.002988,   0.002988,    0.002988,    0.002988,
  0.002988,   0.002988,    0.002988,    0.002988,
  0.002985,   0.002985,    0.002985,    0.002985,
  0.003007,   0.003007,    0.003007,    0.003007,
  0.003013,   0.003013,    0.003013,    0.003013,
  0.002992,   0.002992,    0.002992,    0.002992,
  0.003022,   0.003022,    0.003022,    0.003022,
  0.003101,   0.003101,    0.003101,    0.003101,
  0.003212,   0.003212,    0.003212,    0.003212,
  0.003423,   0.003423,    0.003423,    0.003423,
  0.0036,     0.0036,      0.0036,      0.0036,
  0.003721,   0.003721,    0.003721,    0.003721,
  0.003982,   0.003982,    0.003982,    0.003982,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004448,   0.004448,    0.004448,    0.004448,
  0.004656,   0.004656,    0.004656,    0.004656,
  0.004688,   0.004688,    0.004688,    0.004688,
  0.004684,   0.004684,    0.004684,    0.004684,
  0.004792,   0.004792,    0.004792,    0.004792,
  0.004949,   0.004949,    0.004949,    0.004949,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005154,   0.005154,    0.005154,    0.005154,
  0.005218,   0.005218,    0.005218,    0.005218,
  0.005266,   0.005266,    0.005266,    0.005266,
  0.005299,   0.005299,    0.005299,    0.005299,
  0.005331,   0.005331,    0.005331,    0.005331,
  0.005397,   0.005397,    0.005397,    0.005397,
  0.0055,     0.0055,      0.0055,      0.0055,
  0.005556,   0.005556,    0.005556,    0.005556,
  0.005612,   0.005612,    0.005612,    0.005612,
  0.005686,   0.005686,    0.005686,    0.005686,
  0.005708,   0.005708,    0.005708,    0.005708,
  0.005708,   0.005708,    0.005708,    0.005708,
  0.005668,   0.005668,    0.005668,    0.005668,
  0.005633,   0.005633,    0.005633,    0.005633,
  0.005677,   0.005677,    0.005677,    0.005677,
  0.005745,   0.005745,    0.005745,    0.005745,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.005737,   0.005737,    0.005737,    0.005737,
  0.005732,   0.005732,    0.005732,    0.005732,
  0.005769,   0.005769,    0.005769,    0.005769,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.005861,   0.005861,    0.005861,    0.005861,
  0.005949,   0.005949,    0.005949,    0.005949,
  0.006038,   0.006038,    0.006038,    0.006038,
  0.006127,   0.006127,    0.006127,    0.006127,
  0.006133,   0.006133,    0.006133,    0.006133,
  0.006133,   0.006133,    0.006133,    0.006133,
  0.006184,   0.006184,    0.006184,    0.006184,
  0.006223,   0.006223,    0.006223,    0.006223,
  0.006235,   0.006235,    0.006235,    0.006235,
  0.006209,   0.006209,    0.006209,    0.006209,
  0.006209,   0.006209,    0.006209,    0.006209,
  0.006216,   0.006216,    0.006216,    0.006216,
  0.006191,   0.006191,    0.006191,    0.006191,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.006153,   0.006153,    0.006153,    0.006153,
  0.006196,   0.006196,    0.006196,    0.006196,
  0.006209,   0.006209,    0.006209,    0.006209,
  0.006151,   0.006151,    0.006151,    0.006151,
  0.006126,   0.006126,    0.006126,    0.006126,
  0.006126,   0.006126,    0.006126,    0.006126,
  0.006132,   0.006132,    0.006132,    0.006132,
  0.006177,   0.006177,    0.006177,    0.006177,
  0.006179,   0.006179,    0.006179,    0.006179,
  0.006143,   0.006143,    0.006143,    0.006143,
  0.006117,   0.006117,    0.006117,    0.006117,
  0.00609,    0.00609,     0.00609,     0.00609,
  0.00612,    0.00612,     0.00612,     0.00612,
  0.006097,   0.006097,    0.006097,    0.006097,
  0.006003,   0.006003,    0.006003,    0.006003,
  0.005971,   0.005971,    0.005971,    0.005971,
  0.005919,   0.005919,    0.005919,    0.005919,
  0.005879,   0.005879,    0.005879,    0.005879,
  0.005893,   0.005893,    0.005893,    0.005893,
  0.005907,   0.005907,    0.005907,    0.005907,
  0.005931,   0.005931,    0.005931,    0.005931,
  0.005931,   0.005931,    0.005931,    0.005931,
  0.005919,   0.005919,    0.005919,    0.005919,
  0.006006,   0.006006,    0.006006,    0.006006,
  0.006172,   0.006172,    0.006172,    0.006172,
  0.006271,   0.006271,    0.006271,    0.006271,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006334,   0.006334,    0.006334,    0.006334,
  0.006391,   0.006391,    0.006391,    0.006391,
  0.00648,    0.00648,     0.00648,     0.00648,
  0.006538,   0.006538,    0.006538,    0.006538,
  0.006596,   0.006596,    0.006596,    0.006596,
  0.006675,   0.006675,    0.006675,    0.006675,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006775,   0.006775,    0.006775,    0.006775,
  0.006795,   0.006795,    0.006795,    0.006795,
  0.006795,   0.006795,    0.006795,    0.006795,
  0.006815,   0.006815,    0.006815,    0.006815,
  0.006855,   0.006855,    0.006855,    0.006855,
  0.006937,   0.006937,    0.006937,    0.006937,
  0.007019,   0.007019,    0.007019,    0.007019,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.007144,   0.007144,    0.007144,    0.007144,
  0.007186,   0.007186,    0.007186,    0.007186,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007186,   0.007186,    0.007186,    0.007186,
  0.007154,   0.007154,    0.007154,    0.007154,
  0.007112,   0.007112,    0.007112,    0.007112,
  0.007028,   0.007028,    0.007028,    0.007028,
  0.006944,   0.006944,    0.006944,    0.006944,
  0.006892,   0.006892,    0.006892,    0.006892,
  0.006851,   0.006851,    0.006851,    0.006851,
  0.006841,   0.006841,    0.006841,    0.006841,
  0.00682,    0.00682,     0.00682,     0.00682,
  0.006829,   0.006829,    0.006829,    0.006829,
  0.006924,   0.006924,    0.006924,    0.006924,
  0.006987,   0.006987,    0.006987,    0.006987,
  0.006998,   0.006998,    0.006998,    0.006998,
  0.007019,   0.007019,    0.007019,    0.007019,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007271,   0.007271,    0.007271,    0.007271,
  0.007378,   0.007378,    0.007378,    0.007378,
  0.007465,   0.007465,    0.007465,    0.007465,
  0.007575,   0.007575,    0.007575,    0.007575,
  0.007731,   0.007731,    0.007731,    0.007731,
  0.007867,   0.007867,    0.007867,    0.007867,
  0.007896,   0.007896,    0.007896,    0.007896,
  0.007816,   0.007816,    0.007816,    0.007816,
  0.007621,   0.007621,    0.007621,    0.007621,
  0.00743,    0.00743,     0.00743,     0.00743,
  0.007326,   0.007326,    0.007326,    0.007326,
  0.007219,   0.007219,    0.007219,    0.007219,
  0.007106,   0.007106,    0.007106,    0.007106,
  0.006971,   0.006971,    0.006971,    0.006971,
  0.006885,   0.006885,    0.006885,    0.006885,
  0.006885,   0.006885,    0.006885,    0.006885,
  0.006885,   0.006885,    0.006885,    0.006885,
  0.006898,   0.006898,    0.006898,    0.006898,
  0.006871,   0.006871,    0.006871,    0.006871,
  0.006871,   0.006871,    0.006871,    0.006871,
  0.006898,   0.006898,    0.006898,    0.006898,
  0.0068,     0.0068,      0.0068,      0.0068,
  0.006806,   0.006806,    0.006806,    0.006806,
  0.006908,   0.006908,    0.006908,    0.006908,
  0.006823,   0.006823,    0.006823,    0.006823,
  0.006612,   0.006612,    0.006612,    0.006612,
  0.006506,   0.006506,    0.006506,    0.006506,
  0.006652,   0.006652,    0.006652,    0.006652,
  0.006798,   0.006798,    0.006798,    0.006798,
  0.006839,   0.006839,    0.006839,    0.006839,
  0.006923,   0.006923,    0.006923,    0.006923,
  0.006986,   0.006986,    0.006986,    0.006986,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007197,   0.007197,    0.007197,    0.007197,
  0.007145,   0.007145,    0.007145,    0.007145,
  0.007103,   0.007103,    0.007103,    0.007103,
  0.007102,   0.007102,    0.007102,    0.007102,
  0.007091,   0.007091,    0.007091,    0.007091,
  0.007081,   0.007081,    0.007081,    0.007081,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.00706,    0.00706,     0.00706,     0.00706,
  0.007165,   0.007165,    0.007165,    0.007165,
  0.007335,   0.007335,    0.007335,    0.007335,
  0.007554,   0.007554,    0.007554,    0.007554,
  0.007736,   0.007736,    0.007736,    0.007736,
  0.007707,   0.007707,    0.007707,    0.007707,
  0.007556,   0.007556,    0.007556,    0.007556,
  0.007405,   0.007405,    0.007405,    0.007405,
  0.007358,   0.007358,    0.007358,    0.007358,
  0.007303,   0.007303,    0.007303,    0.007303,
  0.007201,   0.007201,    0.007201,    0.007201,
  0.007194,   0.007194,    0.007194,    0.007194,
  0.00714,    0.00714,     0.00714,     0.00714,
  0.007054,   0.007054,    0.007054,    0.007054,
  0.007016,   0.007016,    0.007016,    0.007016,
  0.00702,    0.00702,     0.00702,     0.00702,
  0.006975,   0.006975,    0.006975,    0.006975,
  0.006912,   0.006912,    0.006912,    0.006912,
  0.006898,   0.006898,    0.006898,    0.006898,
  0.006882,   0.006882,    0.006882,    0.006882,
  0.006918,   0.006918,    0.006918,    0.006918,
  0.006977,   0.006977,    0.006977,    0.006977,
  0.006914,   0.006914,    0.006914,    0.006914,
  0.006809,   0.006809,    0.006809,    0.006809,
  0.006767,   0.006767,    0.006767,    0.006767,
  0.006745,   0.006745,    0.006745,    0.006745,
  0.006693,   0.006693,    0.006693,    0.006693,
  0.006536,   0.006536,    0.006536,    0.006536,
  0.006361,   0.006361,    0.006361,    0.006361,
  0.006337,   0.006337,    0.006337,    0.006337,
  0.006376,   0.006376,    0.006376,    0.006376,
  0.006368,   0.006368,    0.006368,    0.006368,
  0.006368,   0.006368,    0.006368,    0.006368,
  0.006412,   0.006412,    0.006412,    0.006412,
  0.006468,   0.006468,    0.006468,    0.006468,
  0.006423,   0.006423,    0.006423,    0.006423,
  0.00629,    0.00629,     0.00629,     0.00629,
  0.006197,   0.006197,    0.006197,    0.006197,
  0.006178,   0.006178,    0.006178,    0.006178,
  0.006253,   0.006253,    0.006253,    0.006253,
  0.006346,   0.006346,    0.006346,    0.006346,
  0.006384,   0.006384,    0.006384,    0.006384,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006197,   0.006197,    0.006197,    0.006197,
  0.00616,    0.00616,     0.00616,     0.00616,
  0.006068,   0.006068,    0.006068,    0.006068,
  0.00596,    0.00596,     0.00596,     0.00596,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005942,   0.005942,    0.005942,    0.005942,
  0.005982,   0.005982,    0.005982,    0.005982,
  0.006028,   0.006028,    0.006028,    0.006028,
  0.006047,   0.006047,    0.006047,    0.006047,
  0.006023,   0.006023,    0.006023,    0.006023,
  0.006023,   0.006023,    0.006023,    0.006023,
  0.006015,   0.006015,    0.006015,    0.006015,
  0.005945,   0.005945,    0.005945,    0.005945,
  0.005869,   0.005869,    0.005869,    0.005869,
  0.005824,   0.005824,    0.005824,    0.005824,
  0.005793,   0.005793,    0.005793,    0.005793,
  0.005813,   0.005813,    0.005813,    0.005813,
  0.005875,   0.005875,    0.005875,    0.005875,
  0.005861,   0.005861,    0.005861,    0.005861,
  0.005843,   0.005843,    0.005843,    0.005843,
  0.005861,   0.005861,    0.005861,    0.005861,
  0.005826,   0.005826,    0.005826,    0.005826,
  0.005755,   0.005755,    0.005755,    0.005755,
  0.005608,   0.005608,    0.005608,    0.005608,
  0.005433,   0.005433,    0.005433,    0.005433,
  0.005325,   0.005325,    0.005325,    0.005325,
  0.005199,   0.005199,    0.005199,    0.005199,
  0.005081,   0.005081,    0.005081,    0.005081,
  0.005072,   0.005072,    0.005072,    0.005072,
  0.005082,   0.005082,    0.005082,    0.005082,
  0.005055,   0.005055,    0.005055,    0.005055,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004715,   0.004715,    0.004715,    0.004715,
  0.004536,   0.004536,    0.004536,    0.004536,
  0.004483,   0.004483,    0.004483,    0.004483,
  0.004448,   0.004448,    0.004448,    0.004448,
  0.004433,   0.004433,    0.004433,    0.004433,
  0.004415,   0.004415,    0.004415,    0.004415,
  0.004384,   0.004384,    0.004384,    0.004384,
  0.004371,   0.004371,    0.004371,    0.004371,
  0.004389,   0.004389,    0.004389,    0.004389,
  0.004437,   0.004437,    0.004437,    0.004437,
  0.004471,   0.004471,    0.004471,    0.004471,
  0.004489,   0.004489,    0.004489,    0.004489,
  0.00455,    0.00455,     0.00455,     0.00455,
  0.004671,   0.004671,    0.004671,    0.004671,
  0.004794,   0.004794,    0.004794,    0.004794,
  0.004841,   0.004841,    0.004841,    0.004841,
  0.004796,   0.004796,    0.004796,    0.004796,
  0.004706,   0.004706,    0.004706,    0.004706,
  0.004661,   0.004661,    0.004661,    0.004661,
  0.004661,   0.004661,    0.004661,    0.004661,
  0.00472,    0.00472,     0.00472,     0.00472,
  0.004824,   0.004824,    0.004824,    0.004824,
  0.004986,   0.004986,    0.004986,    0.004986,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005331,   0.005331,    0.005331,    0.005331,
  0.005377,   0.005377,    0.005377,    0.005377,
  0.005357,   0.005357,    0.005357,    0.005357,
  0.005401,   0.005401,    0.005401,    0.005401,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005578,   0.005578,    0.005578,    0.005578,
  0.005745,   0.005745,    0.005745,    0.005745,
  0.005874,   0.005874,    0.005874,    0.005874,
  0.005924,   0.005924,    0.005924,    0.005924,
  0.005979,   0.005979,    0.005979,    0.005979,
  0.005984,   0.005984,    0.005984,    0.005984,
  0.005971,   0.005971,    0.005971,    0.005971,
  0.00602,    0.00602,     0.00602,     0.00602,
  0.006052,   0.006052,    0.006052,    0.006052,
  0.006034,   0.006034,    0.006034,    0.006034,
  0.006015,   0.006015,    0.006015,    0.006015,
  0.006028,   0.006028,    0.006028,    0.006028,
  0.006005,   0.006005,    0.006005,    0.006005,
  0.005964,   0.005964,    0.005964,    0.005964,
  0.005907,   0.005907,    0.005907,    0.005907,
  0.005818,   0.005818,    0.005818,    0.005818,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005679,   0.005679,    0.005679,    0.005679,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.00556,    0.00556,     0.00556,     0.00556,
  0.005494,   0.005494,    0.005494,    0.005494,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005394,   0.005394,    0.005394,    0.005394,
  0.005411,   0.005411,    0.005411,    0.005411,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.004968,   0.004968,    0.004968,    0.004968,
  0.004877,   0.004877,    0.004877,    0.004877,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004802,   0.004802,    0.004802,    0.004802,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.005156,   0.005156,    0.005156,    0.005156,
  0.005151,   0.005151,    0.005151,    0.005151,
  0.004902,   0.004902,    0.004902,    0.004902,
  0.004723,   0.004723,    0.004723,    0.004723,
  0.004651,   0.004651,    0.004651,    0.004651,
  0.004623,   0.004623,    0.004623,    0.004623,
  0.00457,    0.00457,     0.00457,     0.00457,
  0.00445,    0.00445,     0.00445,     0.00445,
  0.004457,   0.004457,    0.004457,    0.004457,
  0.004531,   0.004531,    0.004531,    0.004531,
  0.00474,    0.00474,     0.00474,     0.00474,
  0.004871,   0.004871,    0.004871,    0.004871,
  0.004776,   0.004776,    0.004776,    0.004776,
  0.004666,   0.004666,    0.004666,    0.004666,
  0.004526,   0.004526,    0.004526,    0.004526,
  0.004385,   0.004385,    0.004385,    0.004385,
  0.004307,   0.004307,    0.004307,    0.004307,
  0.004323,   0.004323,    0.004323,    0.004323,
  0.004323,   0.004323,    0.004323,    0.004323,
  0.004292,   0.004292,    0.004292,    0.004292,
  0.004293,   0.004293,    0.004293,    0.004293,
  0.004248,   0.004248,    0.004248,    0.004248,
  0.004128,   0.004128,    0.004128,    0.004128,
  0.003998,   0.003998,    0.003998,    0.003998,
  0.003934,   0.003934,    0.003934,    0.003934,
  0.0039,     0.0039,      0.0039,      0.0039,
  0.003863,   0.003863,    0.003863,    0.003863,
  0.003845,   0.003845,    0.003845,    0.003845,
  0.003707,   0.003707,    0.003707,    0.003707,
  0.00359,    0.00359,     0.00359,     0.00359,
  0.003603,   0.003603,    0.003603,    0.003603,
  0.003618,   0.003618,    0.003618,    0.003618,
  0.003613,   0.003613,    0.003613,    0.003613,
  0.003612,   0.003612,    0.003612,    0.003612,
  0.003688,   0.003688,    0.003688,    0.003688,
  0.003809,   0.003809,    0.003809,    0.003809,
  0.003945,   0.003945,    0.003945,    0.003945,
  0.004052,   0.004052,    0.004052,    0.004052,
  0.004085,   0.004085,    0.004085,    0.004085,
  0.004018,   0.004018,    0.004018,    0.004018,
  0.003846,   0.003846,    0.003846,    0.003846,
  0.003679,   0.003679,    0.003679,    0.003679,
  0.00349,    0.00349,     0.00349,     0.00349,
  0.003239,   0.003239,    0.003239,    0.003239,
  0.003087,   0.003087,    0.003087,    0.003087,
  0.003113,   0.003113,    0.003113,    0.003113,
  0.003184,   0.003184,    0.003184,    0.003184,
  0.003179,   0.003179,    0.003179,    0.003179,
  0.003148,   0.003148,    0.003148,    0.003148,
  0.003161,   0.003161,    0.003161,    0.003161,
  0.003202,   0.003202,    0.003202,    0.003202,
  0.003193,   0.003193,    0.003193,    0.003193,
  0.003139,   0.003139,    0.003139,    0.003139,
  0.00309,    0.00309,     0.00309,     0.00309,
  0.003059,   0.003059,    0.003059,    0.003059,
  0.003045,   0.003045,    0.003045,    0.003045,
  0.003049,   0.003049,    0.003049,    0.003049,
  0.003053,   0.003053,    0.003053,    0.003053,
  0.002999,   0.002999,    0.002999,    0.002999,
  0.00295,    0.00295,     0.00295,     0.00295,
  0.002929,   0.002929,    0.002929,    0.002929,
  0.002921,   0.002921,    0.002921,    0.002921,
  0.002933,   0.002933,    0.002933,    0.002933,
  0.002957,   0.002957,    0.002957,    0.002957,
  0.002963,   0.002963,    0.002963,    0.002963,
  0.002913,   0.002913,    0.002913,    0.002913,
  0.00287,    0.00287,     0.00287,     0.00287,
  0.002859,   0.002859,    0.002859,    0.002859,
  0.002843,   0.002843,    0.002843,    0.002843,
  0.00285,    0.00285,     0.00285,     0.00285,
  0.002854,   0.002854,    0.002854,    0.002854,
  0.002835,   0.002835,    0.002835,    0.002835,
  0.00283,    0.00283,     0.00283,     0.00283,
  0.002825,   0.002825,    0.002825,    0.002825,
  0.002791,   0.002791,    0.002791,    0.002791,
  0.002778,   0.002778,    0.002778,    0.002778,
  0.002788,   0.002788,    0.002788,    0.002788,
  0.002756,   0.002756,    0.002756,    0.002756,
  0.002703,   0.002703,    0.002703,    0.002703,
  0.002672,   0.002672,    0.002672,    0.002672,
  0.002682,   0.002682,    0.002682,    0.002682,
  0.002693,   0.002693,    0.002693,    0.002693,
  0.002693,   0.002693,    0.002693,    0.002693,
  0.002704,   0.002704,    0.002704,    0.002704,
  0.002725,   0.002725,    0.002725,    0.002725,
  0.002705,   0.002705,    0.002705,    0.002705,
  0.002705,   0.002705,    0.002705,    0.002705,
  0.002683,   0.002683,    0.002683,    0.002683,
  0.002619,   0.002619,    0.002619,    0.002619,
  0.002598,   0.002598,    0.002598,    0.002598,
  0.002556,   0.002556,    0.002556,    0.002556,
  0.002504,   0.002504,    0.002504,    0.002504,
  0.002462,   0.002462,    0.002462,    0.002462,
  0.002431,   0.002431,    0.002431,    0.002431,
  0.00242,    0.00242,     0.00242,     0.00242,
  0.00241,    0.00241,     0.00241,     0.00241,
  0.00234,    0.00234,     0.00234,     0.00234,
  0.002231,   0.002231,    0.002231,    0.002231,
  0.002173,   0.002173,    0.002173,    0.002173,
  0.002141,   0.002141,    0.002141,    0.002141,
  0.002117,   0.002117,    0.002117,    0.002117,
  0.002136,   0.002136,    0.002136,    0.002136,
  0.002139,   0.002139,    0.002139,    0.002139,
  0.002119,   0.002119,    0.002119,    0.002119,
  0.002119,   0.002119,    0.002119,    0.002119,
  0.002132,   0.002132,    0.002132,    0.002132,
  0.002125,   0.002125,    0.002125,    0.002125,
  0.00211,    0.00211,     0.00211,     0.00211,
  0.002087,   0.002087,    0.002087,    0.002087,
  0.00205,    0.00205,     0.00205,     0.00205,
  0.002046,   0.002046,    0.002046,    0.002046,
  0.002065,   0.002065,    0.002065,    0.002065,
  0.002079,   0.002079,    0.002079,    0.002079,
  0.002093,   0.002093,    0.002093,    0.002093,
  0.002098,   0.002098,    0.002098,    0.002098,
  0.002081,   0.002081,    0.002081,    0.002081,
  0.002064,   0.002064,    0.002064,    0.002064,
  0.002087,   0.002087,    0.002087,    0.002087,
  0.002119,   0.002119,    0.002119,    0.002119,
  0.002102,   0.002102,    0.002102,    0.002102,
  0.0021,     0.0021,      0.0021,      0.0021,
  0.002106,   0.002106,    0.002106,    0.002106,
  0.002098,   0.002098,    0.002098,    0.002098,
  0.002082,   0.002082,    0.002082,    0.002082,
  0.002057,   0.002057,    0.002057,    0.002057,
  0.002041,   0.002041,    0.002041,    0.002041,
  0.002025,   0.002025,    0.002025,    0.002025,
  0.001985,   0.001985,    0.001985,    0.001985,
  0.001954,   0.001954,    0.001954,    0.001954,
  0.001962,   0.001962,    0.001962,    0.001962,
  0.001938,   0.001938,    0.001938,    0.001938,
  0.001907,   0.001907,    0.001907,    0.001907,
  0.001899,   0.001899,    0.001899,    0.001899,
  0.001883,   0.001883,    0.001883,    0.001883,
  0.001875,   0.001875,    0.001875,    0.001875,
  0.001867,   0.001867,    0.001867,    0.001867,
  0.001859,   0.001859,    0.001859,    0.001859,
  0.001867,   0.001867,    0.001867,    0.001867,
  0.001875,   0.001875,    0.001875,    0.001875,
  0.001883,   0.001883,    0.001883,    0.001883,
  0.001891,   0.001891,    0.001891,    0.001891,
  0.001899,   0.001899,    0.001899,    0.001899,
  0.0019,     0.0019,      0.0019,      0.0019,
  0.001926,   0.001926,    0.001926,    0.001926,
  0.001961,   0.001961,    0.001961,    0.001961,
  0.001985,   0.001985,    0.001985,    0.001985,
  0.002019,   0.002019,    0.002019,    0.002019,
  0.002051,   0.002051,    0.002051,    0.002051,
  0.002075,   0.002075,    0.002075,    0.002075,
  0.002098,   0.002098,    0.002098,    0.002098,
  0.002132,   0.002132,    0.002132,    0.002132,
  0.002181,   0.002181,    0.002181,    0.002181,
  0.002242,   0.002242,    0.002242,    0.002242,
  0.002283,   0.002283,    0.002283,    0.002283,
  0.002336,   0.002336,    0.002336,    0.002336,
  0.002368,   0.002368,    0.002368,    0.002368,
  0.00239,    0.00239,     0.00239,     0.00239,
  0.002411,   0.002411,    0.002411,    0.002411,
  0.002412,   0.002412,    0.002412,    0.002412,
  0.002423,   0.002423,    0.002423,    0.002423,
  0.002455,   0.002455,    0.002455,    0.002455,
  0.002507,   0.002507,    0.002507,    0.002507,
  0.002528,   0.002528,    0.002528,    0.002528,
  0.002507,   0.002507,    0.002507,    0.002507,
  0.002486,   0.002486,    0.002486,    0.002486,
  0.002486,   0.002486,    0.002486,    0.002486,
  0.002497,   0.002497,    0.002497,    0.002497,
  0.00252,    0.00252,     0.00252,     0.00252,
  0.002531,   0.002531,    0.002531,    0.002531,
  0.002573,   0.002573,    0.002573,    0.002573,
  0.002627,   0.002627,    0.002627,    0.002627,
  0.00265,    0.00265,     0.00265,     0.00265,
  0.002684,   0.002684,    0.002684,    0.002684,
  0.002741,   0.002741,    0.002741,    0.002741,
  0.002791,   0.002791,    0.002791,    0.002791,
  0.002831,   0.002831,    0.002831,    0.002831,
  0.002879,   0.002879,    0.002879,    0.002879,
  0.002959,   0.002959,    0.002959,    0.002959,
  0.003027,   0.003027,    0.003027,    0.003027,
  0.003059,   0.003059,    0.003059,    0.003059,
  0.003109,   0.003109,    0.003109,    0.003109,
  0.003159,   0.003159,    0.003159,    0.003159,
  0.003223,   0.003223,    0.003223,    0.003223,
  0.003312,   0.003312,    0.003312,    0.003312,
  0.003375,   0.003375,    0.003375,    0.003375,
  0.003381,   0.003381,    0.003381,    0.003381,
  0.003394,   0.003394,    0.003394,    0.003394,
  0.00345,    0.00345,     0.00345,     0.00345,
  0.003463,   0.003463,    0.003463,    0.003463,
  0.003481,   0.003481,    0.003481,    0.003481,
  0.003564,   0.003564,    0.003564,    0.003564,
  0.00362,    0.00362,     0.00362,     0.00362,
  0.003671,   0.003671,    0.003671,    0.003671,
  0.00371,    0.00371,     0.00371,     0.00371,
  0.00369,    0.00369,     0.00369,     0.00369,
  0.003689,   0.003689,    0.003689,    0.003689,
  0.00372,    0.00372,     0.00372,     0.00372,
  0.003799,   0.003799,    0.003799,    0.003799,
  0.003894,   0.003894,    0.003894,    0.003894,
  0.003895,   0.003895,    0.003895,    0.003895,
  0.003849,   0.003849,    0.003849,    0.003849,
  0.00385,    0.00385,     0.00385,     0.00385,
  0.003854,   0.003854,    0.003854,    0.003854,
  0.003872,   0.003872,    0.003872,    0.003872,
  0.003992,   0.003992,    0.003992,    0.003992,
  0.004177,   0.004177,    0.004177,    0.004177,
  0.004256,   0.004256,    0.004256,    0.004256,
  0.004209,   0.004209,    0.004209,    0.004209,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.00415,    0.00415,     0.00415,     0.00415,
  0.004167,   0.004167,    0.004167,    0.004167,
  0.004263,   0.004263,    0.004263,    0.004263,
  0.00434,    0.00434,     0.00434,     0.00434,
  0.004352,   0.004352,    0.004352,    0.004352,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004256,   0.004256,    0.004256,    0.004256,
  0.004209,   0.004209,    0.004209,    0.004209,
  0.004273,   0.004273,    0.004273,    0.004273,
  0.004369,   0.004369,    0.004369,    0.004369,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004462,   0.004462,    0.004462,    0.004462,
  0.004446,   0.004446,    0.004446,    0.004446,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004508,   0.004508,    0.004508,    0.004508,
  0.004635,   0.004635,    0.004635,    0.004635,
  0.00478,    0.00478,     0.00478,     0.00478,
  0.004875,   0.004875,    0.004875,    0.004875,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004983,   0.004983,    0.004983,    0.004983,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005346,   0.005346,    0.005346,    0.005346,
  0.005414,   0.005414,    0.005414,    0.005414,
  0.005466,   0.005466,    0.005466,    0.005466,
  0.0055,     0.0055,      0.0055,      0.0055,
  0.005439,   0.005439,    0.005439,    0.005439,
  0.005347,   0.005347,    0.005347,    0.005347,
  0.005287,   0.005287,    0.005287,    0.005287,
  0.005276,   0.005276,    0.005276,    0.005276,
  0.00534,    0.00534,     0.00534,     0.00534,
  0.005468,   0.005468,    0.005468,    0.005468,
  0.005515,   0.005515,    0.005515,    0.005515,
  0.005547,   0.005547,    0.005547,    0.005547,
  0.005572,   0.005572,    0.005572,    0.005572,
  0.005565,   0.005565,    0.005565,    0.005565,
  0.005669,   0.005669,    0.005669,    0.005669,
  0.005845,   0.005845,    0.005845,    0.005845,
  0.006073,   0.006073,    0.006073,    0.006073,
  0.006254,   0.006254,    0.006254,    0.006254,
  0.006073,   0.006073,    0.006073,    0.006073,
  0.005755,   0.005755,    0.005755,    0.005755,
  0.005621,   0.005621,    0.005621,    0.005621,
  0.005553,   0.005553,    0.005553,    0.005553,
  0.005548,   0.005548,    0.005548,    0.005548,
  0.005599,   0.005599,    0.005599,    0.005599,
  0.005664,   0.005664,    0.005664,    0.005664,
  0.005719,   0.005719,    0.005719,    0.005719,
  0.005737,   0.005737,    0.005737,    0.005737,
  0.005719,   0.005719,    0.005719,    0.005719,
  0.005669,   0.005669,    0.005669,    0.005669,
  0.005619,   0.005619,    0.005619,    0.005619,
  0.005596,   0.005596,    0.005596,    0.005596,
  0.005533,   0.005533,    0.005533,    0.005533,
  0.005454,   0.005454,    0.005454,    0.005454,
  0.005382,   0.005382,    0.005382,    0.005382,
  0.005296,   0.005296,    0.005296,    0.005296,
  0.005227,   0.005227,    0.005227,    0.005227,
  0.005158,   0.005158,    0.005158,    0.005158,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005012,   0.005012,    0.005012,    0.005012,
  0.004936,   0.004936,    0.004936,    0.004936,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004176,   0.004176,    0.004176,    0.004176,
  0.004163,   0.004163,    0.004163,    0.004163,
  0.004256,   0.004256,    0.004256,    0.004256,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004529,   0.004529,    0.004529,    0.004529,
  0.004642,   0.004642,    0.004642,    0.004642,
  0.004759,   0.004759,    0.004759,    0.004759,
  0.004953,   0.004953,    0.004953,    0.004953,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005187,   0.005187,    0.005187,    0.005187,
  0.005221,   0.005221,    0.005221,    0.005221,
  0.005189,   0.005189,    0.005189,    0.005189,
  0.005124,   0.005124,    0.005124,    0.005124,
  0.004982,   0.004982,    0.004982,    0.004982,
  0.004787,   0.004787,    0.004787,    0.004787,
  0.004628,   0.004628,    0.004628,    0.004628,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004515,   0.004515,    0.004515,    0.004515,
  0.004628,   0.004628,    0.004628,    0.004628,
  0.004656,   0.004656,    0.004656,    0.004656,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004657,   0.004657,    0.004657,    0.004657,
  0.004543,   0.004543,    0.004543,    0.004543,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004473,   0.004473,    0.004473,    0.004473,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004309,   0.004309,    0.004309,    0.004309,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004472,   0.004472,    0.004472,    0.004472,
  0.004472,   0.004472,    0.004472,    0.004472,
  0.004472,   0.004472,    0.004472,    0.004472,
  0.004472,   0.004472,    0.004472,    0.004472,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004473,   0.004473,    0.004473,    0.004473,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004472,   0.004472,    0.004472,    0.004472,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004486,   0.004486,    0.004486,    0.004486,
  0.004472,   0.004472,    0.004472,    0.004472,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004445,   0.004445,    0.004445,    0.004445,
  0.004417,   0.004417,    0.004417,    0.004417,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004336,   0.004336,    0.004336,    0.004336,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.00439,    0.00439,     0.00439,     0.00439,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004363,   0.004363,    0.004363,    0.004363,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004335,   0.004335,    0.004335,    0.004335,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004308,   0.004308,    0.004308,    0.004308,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004308,   0.004308,    0.004308,    0.004308,
  0.004308,   0.004308,    0.004308,    0.004308,
  0.004308,   0.004308,    0.004308,    0.004308,
  0.004308,   0.004308,    0.004308,    0.004308,
  0.004308,   0.004308,    0.004308,    0.004308,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004255,   0.004255,    0.004255,    0.004255,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004202,   0.004202,    0.004202,    0.004202,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004176,   0.004176,    0.004176,    0.004176,
  0.004176,   0.004176,    0.004176,    0.004176,
  0.004189,   0.004189,    0.004189,    0.004189,
  0.004215,   0.004215,    0.004215,    0.004215,
  0.004228,   0.004228,    0.004228,    0.004228,
  0.004242,   0.004242,    0.004242,    0.004242,
  0.004268,   0.004268,    0.004268,    0.004268,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004431,   0.004431,    0.004431,    0.004431,
  0.004473,   0.004473,    0.004473,    0.004473,
  0.004514,   0.004514,    0.004514,    0.004514,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004528,   0.004528,    0.004528,    0.004528,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004542,   0.004542,    0.004542,    0.004542,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004671,   0.004671,    0.004671,    0.004671,
  0.004744,   0.004744,    0.004744,    0.004744,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.005014,   0.005014,    0.005014,    0.005014,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005265,   0.005265,    0.005265,    0.005265,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005427,   0.005427,    0.005427,    0.005427,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005477,   0.005477,    0.005477,    0.005477,
  0.005493,   0.005493,    0.005493,    0.005493,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.00556,    0.00556,     0.00556,     0.00556,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005697,   0.005697,    0.005697,    0.005697,
  0.005801,   0.005801,    0.005801,    0.005801,
  0.005907,   0.005907,    0.005907,    0.005907,
  0.00605,    0.00605,     0.00605,     0.00605,
  0.006253,   0.006253,    0.006253,    0.006253,
  0.006481,   0.006481,    0.006481,    0.006481,
  0.006656,   0.006656,    0.006656,    0.006656,
  0.006775,   0.006775,    0.006775,    0.006775,
  0.006876,   0.006876,    0.006876,    0.006876,
  0.006999,   0.006999,    0.006999,    0.006999,
  0.007123,   0.007123,    0.007123,    0.007123,
  0.007207,   0.007207,    0.007207,    0.007207,
  0.007249,   0.007249,    0.007249,    0.007249,
  0.007271,   0.007271,    0.007271,    0.007271,
  0.007335,   0.007335,    0.007335,    0.007335,
  0.0074,     0.0074,      0.0074,      0.0074,
  0.007443,   0.007443,    0.007443,    0.007443,
  0.007509,   0.007509,    0.007509,    0.007509,
  0.007575,   0.007575,    0.007575,    0.007575,
  0.007597,   0.007597,    0.007597,    0.007597,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007664,   0.007664,    0.007664,    0.007664,
  0.007708,   0.007708,    0.007708,    0.007708,
  0.007731,   0.007731,    0.007731,    0.007731,
  0.007731,   0.007731,    0.007731,    0.007731,
  0.007753,   0.007753,    0.007753,    0.007753,
  0.007776,   0.007776,    0.007776,    0.007776,
  0.007799,   0.007799,    0.007799,    0.007799,
  0.007844,   0.007844,    0.007844,    0.007844,
  0.007821,   0.007821,    0.007821,    0.007821,
  0.007753,   0.007753,    0.007753,    0.007753,
  0.007686,   0.007686,    0.007686,    0.007686,
  0.007619,   0.007619,    0.007619,    0.007619,
  0.007553,   0.007553,    0.007553,    0.007553,
  0.007465,   0.007465,    0.007465,    0.007465,
  0.007421,   0.007421,    0.007421,    0.007421,
  0.007455,   0.007455,    0.007455,    0.007455,
  0.007471,   0.007471,    0.007471,    0.007471,
  0.00738,    0.00738,     0.00738,     0.00738,
  0.007209,   0.007209,    0.007209,    0.007209,
  0.006985,   0.006985,    0.006985,    0.006985,
  0.006809,   0.006809,    0.006809,    0.006809,
  0.006687,   0.006687,    0.006687,    0.006687,
  0.006381,   0.006381,    0.006381,    0.006381,
  0.00606,    0.00606,     0.00606,     0.00606,
  0.005908,   0.005908,    0.005908,    0.005908,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005821,   0.005821,    0.005821,    0.005821,
  0.005716,   0.005716,    0.005716,    0.005716,
  0.005696,   0.005696,    0.005696,    0.005696,
  0.005783,   0.005783,    0.005783,    0.005783,
  0.005838,   0.005838,    0.005838,    0.005838,
  0.00583,    0.00583,     0.00583,     0.00583,
  0.00581,    0.00581,     0.00581,     0.00581,
  0.005821,   0.005821,    0.005821,    0.005821,
  0.005805,   0.005805,    0.005805,    0.005805,
  0.005797,   0.005797,    0.005797,    0.005797,
  0.005817,   0.005817,    0.005817,    0.005817,
  0.005828,   0.005828,    0.005828,    0.005828,
  0.005821,   0.005821,    0.005821,    0.005821,
  0.005821,   0.005821,    0.005821,    0.005821,
  0.005797,   0.005797,    0.005797,    0.005797,
  0.005762,   0.005762,    0.005762,    0.005762,
  0.005801,   0.005801,    0.005801,    0.005801,
  0.005853,   0.005853,    0.005853,    0.005853,
  0.005913,   0.005913,    0.005913,    0.005913,
  0.005962,   0.005962,    0.005962,    0.005962,
  0.006086,   0.006086,    0.006086,    0.006086,
  0.006274,   0.006274,    0.006274,    0.006274,
  0.006577,   0.006577,    0.006577,    0.006577,
  0.007029,   0.007029,    0.007029,    0.007029,
  0.007382,   0.007382,    0.007382,    0.007382,
  0.007551,   0.007551,    0.007551,    0.007551,
  0.007592,   0.007592,    0.007592,    0.007592,
  0.007644,   0.007644,    0.007644,    0.007644,
  0.007486,   0.007486,    0.007486,    0.007486,
  0.007003,   0.007003,    0.007003,    0.007003,
  0.006632,   0.006632,    0.006632,    0.006632,
  0.006412,   0.006412,    0.006412,    0.006412,
  0.00619,    0.00619,     0.00619,     0.00619,
  0.006042,   0.006042,    0.006042,    0.006042,
  0.005937,   0.005937,    0.005937,    0.005937,
  0.005863,   0.005863,    0.005863,    0.005863,
  0.005884,   0.005884,    0.005884,    0.005884,
  0.005916,   0.005916,    0.005916,    0.005916,
  0.005769,   0.005769,    0.005769,    0.005769,
  0.005632,   0.005632,    0.005632,    0.005632,
  0.00559,    0.00559,     0.00559,     0.00559,
  0.005569,   0.005569,    0.005569,    0.005569,
  0.005538,   0.005538,    0.005538,    0.005538,
  0.005475,   0.005475,    0.005475,    0.005475,
  0.005455,   0.005455,    0.005455,    0.005455,
  0.005445,   0.005445,    0.005445,    0.005445,
  0.005423,   0.005423,    0.005423,    0.005423,
  0.005349,   0.005349,    0.005349,    0.005349,
  0.005266,   0.005266,    0.005266,    0.005266,
  0.005256,   0.005256,    0.005256,    0.005256,
  0.005321,   0.005321,    0.005321,    0.005321,
  0.005321,   0.005321,    0.005321,    0.005321,
  0.005343,   0.005343,    0.005343,    0.005343,
  0.005463,   0.005463,    0.005463,    0.005463,
  0.005475,   0.005475,    0.005475,    0.005475,
  0.005459,   0.005459,    0.005459,    0.005459,
  0.005399,   0.005399,    0.005399,    0.005399,
  0.005392,   0.005392,    0.005392,    0.005392,
  0.005541,   0.005541,    0.005541,    0.005541,
  0.005634,   0.005634,    0.005634,    0.005634,
  0.00561,    0.00561,     0.00561,     0.00561,
  0.005528,   0.005528,    0.005528,    0.005528,
  0.005667,   0.005667,    0.005667,    0.005667,
  0.005832,   0.005832,    0.005832,    0.005832,
  0.005839,   0.005839,    0.005839,    0.005839,
  0.005776,   0.005776,    0.005776,    0.005776,
  0.005648,   0.005648,    0.005648,    0.005648,
  0.005597,   0.005597,    0.005597,    0.005597,
  0.005702,   0.005702,    0.005702,    0.005702,
  0.00582,    0.00582,     0.00582,     0.00582,
  0.00583,    0.00583,     0.00583,     0.00583,
  0.005826,   0.005826,    0.005826,    0.005826,
  0.005826,   0.005826,    0.005826,    0.005826,
  0.005759,   0.005759,    0.005759,    0.005759,
  0.005657,   0.005657,    0.005657,    0.005657,
  0.005602,   0.005602,    0.005602,    0.005602,
  0.005548,   0.005548,    0.005548,    0.005548,
  0.005546,   0.005546,    0.005546,    0.005546,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.00556,    0.00556,     0.00556,     0.00556,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005413,   0.005413,    0.005413,    0.005413,
  0.005298,   0.005298,    0.005298,    0.005298,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005249,   0.005249,    0.005249,    0.005249,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005297,   0.005297,    0.005297,    0.005297,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005249,   0.005249,    0.005249,    0.005249,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005249,   0.005249,    0.005249,    0.005249,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005662,   0.005662,    0.005662,    0.005662,
  0.005548,   0.005548,    0.005548,    0.005548,
  0.005531,   0.005531,    0.005531,    0.005531,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005611,   0.005611,    0.005611,    0.005611,
  0.005512,   0.005512,    0.005512,    0.005512,
  0.005479,   0.005479,    0.005479,    0.005479,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005628,   0.005628,    0.005628,    0.005628,
  0.005594,   0.005594,    0.005594,    0.005594,
  0.005577,   0.005577,    0.005577,    0.005577,
  0.00556,    0.00556,     0.00556,     0.00556,
  0.005544,   0.005544,    0.005544,    0.005544,
  0.005527,   0.005527,    0.005527,    0.005527,
  0.00546,    0.00546,     0.00546,     0.00546,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005153,   0.005153,    0.005153,    0.005153,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.004998,   0.004998,    0.004998,    0.004998,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004758,   0.004758,    0.004758,    0.004758,
  0.004729,   0.004729,    0.004729,    0.004729,
  0.004714,   0.004714,    0.004714,    0.004714,
  0.004657,   0.004657,    0.004657,    0.004657,
  0.004585,   0.004585,    0.004585,    0.004585,
  0.004585,   0.004585,    0.004585,    0.004585,
  0.004686,   0.004686,    0.004686,    0.004686,
  0.004817,   0.004817,    0.004817,    0.004817,
  0.004892,   0.004892,    0.004892,    0.004892,
  0.004952,   0.004952,    0.004952,    0.004952,
  0.005076,   0.005076,    0.005076,    0.005076,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005346,   0.005346,    0.005346,    0.005346,
  0.005364,   0.005364,    0.005364,    0.005364,
  0.005334,   0.005334,    0.005334,    0.005334,
  0.005321,   0.005321,    0.005321,    0.005321,
  0.005306,   0.005306,    0.005306,    0.005306,
  0.00529,    0.00529,     0.00529,     0.00529,
  0.005273,   0.005273,    0.005273,    0.005273,
  0.005271,   0.005271,    0.005271,    0.005271,
  0.005222,   0.005222,    0.005222,    0.005222,
  0.005173,   0.005173,    0.005173,    0.005173,
  0.005139,   0.005139,    0.005139,    0.005139,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.005059,   0.005059,    0.005059,    0.005059,
  0.005059,   0.005059,    0.005059,    0.005059,
  0.005091,   0.005091,    0.005091,    0.005091,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005329,   0.005329,    0.005329,    0.005329,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005233,   0.005233,    0.005233,    0.005233,
  0.005201,   0.005201,    0.005201,    0.005201,
  0.005185,   0.005185,    0.005185,    0.005185,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005138,   0.005138,    0.005138,    0.005138,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.00506,    0.00506,     0.00506,     0.00506,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.005028,   0.005028,    0.005028,    0.005028,
  0.005013,   0.005013,    0.005013,    0.005013,
  0.005029,   0.005029,    0.005029,    0.005029,
  0.004953,   0.004953,    0.004953,    0.004953,
  0.004803,   0.004803,    0.004803,    0.004803,
  0.004671,   0.004671,    0.004671,    0.004671,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.0045,     0.0045,      0.0045,      0.0045,
  0.004557,   0.004557,    0.004557,    0.004557,
  0.00473,    0.00473,     0.00473,     0.00473,
  0.004876,   0.004876,    0.004876,    0.004876,
  0.004966,   0.004966,    0.004966,    0.004966,
  0.005077,   0.005077,    0.005077,    0.005077,
  0.005194,   0.005194,    0.005194,    0.005194,
  0.005268,   0.005268,    0.005268,    0.005268,
  0.005227,   0.005227,    0.005227,    0.005227,
  0.005181,   0.005181,    0.005181,    0.005181,
  0.005144,   0.005144,    0.005144,    0.005144,
  0.005136,   0.005136,    0.005136,    0.005136,
  0.005162,   0.005162,    0.005162,    0.005162,
  0.005125,   0.005125,    0.005125,    0.005125,
  0.005075,   0.005075,    0.005075,    0.005075,
  0.005106,   0.005106,    0.005106,    0.005106,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005362,   0.005362,    0.005362,    0.005362,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005378,   0.005378,    0.005378,    0.005378,
  0.005345,   0.005345,    0.005345,    0.005345,
  0.005313,   0.005313,    0.005313,    0.005313,
  0.005281,   0.005281,    0.005281,    0.005281,
  0.005217,   0.005217,    0.005217,    0.005217,
  0.005169,   0.005169,    0.005169,    0.005169,
  0.005122,   0.005122,    0.005122,    0.005122,
  0.005044,   0.005044,    0.005044,    0.005044,
  0.004968,   0.004968,    0.004968,    0.004968,
  0.004937,   0.004937,    0.004937,    0.004937,
  0.004922,   0.004922,    0.004922,    0.004922,
  0.004847,   0.004847,    0.004847,    0.004847,
  0.004773,   0.004773,    0.004773,    0.004773,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004743,   0.004743,    0.004743,    0.004743,
  0.004685,   0.004685,    0.004685,    0.004685,
  0.004613,   0.004613,    0.004613,    0.004613,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004571,   0.004571,    0.004571,    0.004571,
  0.004543,   0.004543,    0.004543,    0.004543,
  0.004459,   0.004459,    0.004459,    0.004459,
  0.004376,   0.004376,    0.004376,    0.004376,
  0.004309,   0.004309,    0.004309,    0.004309,
  0.004282,   0.004282,    0.004282,    0.004282,
  0.004295,   0.004295,    0.004295,    0.004295,
  0.004322,   0.004322,    0.004322,    0.004322,
  0.004349,   0.004349,    0.004349,    0.004349,
  0.004404,   0.004404,    0.004404,    0.004404,
  0.004515,   0.004515,    0.004515,    0.004515,
  0.00465,    0.00465,     0.00465,     0.00465,
  0.004635,   0.004635,    0.004635,    0.004635,
  0.004556,   0.004556,    0.004556,    0.004556,
  0.004543,   0.004543,    0.004543,    0.004543,
  0.004481,   0.004481,    0.004481,    0.004481,
  0.004449,   0.004449,    0.004449,    0.004449,
  0.004466,   0.004466,    0.004466,    0.004466,
  0.004484,   0.004484,    0.004484,    0.004484,
  0.004507,   0.004507,    0.004507,    0.004507,
  0.004483,   0.004483,    0.004483,    0.004483,
  0.004454,   0.004454,    0.004454,    0.004454,
  0.004485,   0.004485,    0.004485,    0.004485,
  0.004517,   0.004517,    0.004517,    0.004517,
  0.00452,    0.00452,     0.00452,     0.00452,
  0.004527,   0.004527,    0.004527,    0.004527,
  0.004566,   0.004566,    0.004566,    0.004566,
  0.004637,   0.004637,    0.004637,    0.004637,
  0.004722,   0.004722,    0.004722,    0.004722,
  0.00479,    0.00479,     0.00479,     0.00479,
  0.004845,   0.004845,    0.004845,    0.004845,
  0.004913,   0.004913,    0.004913,    0.004913,
  0.004944,   0.004944,    0.004944,    0.004944,
  0.004989,   0.004989,    0.004989,    0.004989,
  0.005052,   0.005052,    0.005052,    0.005052,
  0.005089,   0.005089,    0.005089,    0.005089,
  0.005107,   0.005107,    0.005107,    0.005107,
  0.005089,   0.005089,    0.005089,    0.005089,
  0.00507,    0.00507,     0.00507,     0.00507,
  0.005102,   0.005102,    0.005102,    0.005102,
  0.005215,   0.005215,    0.005215,    0.005215,
  0.005359,   0.005359,    0.005359,    0.005359,
  0.005472,   0.005472,    0.005472,    0.005472,
  0.005528,   0.005528,    0.005528,    0.005528,
  0.005553,   0.005553,    0.005553,    0.005553,
  0.005603,   0.005603,    0.005603,    0.005603,
  0.005653,   0.005653,    0.005653,    0.005653,
  0.005647,   0.005647,    0.005647,    0.005647,
  0.005603,   0.005603,    0.005603,    0.005603,
  0.005578,   0.005578,    0.005578,    0.005578,
  0.005546,   0.005546,    0.005546,    0.005546,
  0.005622,   0.005622,    0.005622,    0.005622,
  0.005786,   0.005786,    0.005786,    0.005786,
  0.00595,    0.00595,     0.00595,     0.00595,
  0.006115,   0.006115,    0.006115,    0.006115,
  0.006234,   0.006234,    0.006234,    0.006234,
  0.006309,   0.006309,    0.006309,    0.006309,
  0.006365,   0.006365,    0.006365,    0.006365,
  0.006442,   0.006442,    0.006442,    0.006442,
  0.006538,   0.006538,    0.006538,    0.006538,
  0.006616,   0.006616,    0.006616,    0.006616,
  0.006655,   0.006655,    0.006655,    0.006655,
  0.006695,   0.006695,    0.006695,    0.006695,
  0.006715,   0.006715,    0.006715,    0.006715,
  0.006715,   0.006715,    0.006715,    0.006715,
  0.006735,   0.006735,    0.006735,    0.006735,
  0.006763,   0.006763,    0.006763,    0.006763,
  0.006772,   0.006772,    0.006772,    0.006772,
  0.00674,    0.00674,     0.00674,     0.00674,
  0.006709,   0.006709,    0.006709,    0.006709,
  0.006669,   0.006669,    0.006669,    0.006669,
  0.006589,   0.006589,    0.006589,    0.006589,
  0.00651,    0.00651,     0.00651,     0.00651,
  0.006349,   0.006349,    0.006349,    0.006349,
  0.006183,   0.006183,    0.006183,    0.006183,
  0.006132,   0.006132,    0.006132,    0.006132,
  0.006121,   0.006121,    0.006121,    0.006121,
  0.006078,   0.006078,    0.006078,    0.006078,
  0.006037,   0.006037,    0.006037,    0.006037,
  0.006014,   0.006014,    0.006014,    0.006014,
  0.005946,   0.005946,    0.005946,    0.005946,
  0.005879,   0.005879,    0.005879,    0.005879,
  0.00584,    0.00584,     0.00584,     0.00584,
  0.005783,   0.005783,    0.005783,    0.005783,
  0.005731,   0.005731,    0.005731,    0.005731,
  0.005697, 0.005697, 0.005697,   0.005697 ;

 Wind =
  2.017,   2.017,   2.017,   2.017,
  3.77,    3.77,    3.77,    3.77,
  4.29,    4.29,    4.29,    4.29,
  4.42,    4.42,    4.42,    4.42,
  4.08,    4.08,    4.08,    4.08,
  3.73,    3.73,    3.73,    3.73,
  4,       4,       4,       4,
  4.36,    4.36,    4.36,    4.36,
  4.38,    4.38,    4.38,    4.38,
  3.92,    3.92,    3.92,    3.92,
  4.16,    4.16,    4.16,    4.16,
  4.07,    4.07,    4.07,    4.07,
  4.47,    4.47,    4.47,    4.47,
  4.2,     4.2,     4.2,     4.2,
  3.95,    3.95,    3.95,    3.95,
  3.99,    3.99,    3.99,    3.99,
  3.74,    3.74,    3.74,    3.74,
  3.61,    3.61,    3.61,    3.61,
  3.01,    3.01,    3.01,    3.01,
  3.14,    3.14,    3.14,    3.14,
  2.89,    2.89,    2.89,    2.89,
  3.6,     3.6,     3.6,     3.6,
  3.24,    3.24,    3.24,    3.24,
  3.14,    3.14,    3.14,    3.14,
  3.29,    3.29,    3.29,    3.29,
  4,       4,       4,       4,
  3.09,    3.09,    3.09,    3.09,
  3.08,    3.08,    3.08,    3.08,
  3.86,    3.86,    3.86,    3.86,
  3.49,    3.49,    3.49,    3.49,
  3.36,    3.36,    3.36,    3.36,
  3.19,    3.19,    3.19,    3.19,
  3.16,    3.16,    3.16,    3.16,
  2.15,    2.15,    2.15,    2.15,
  2.16,    2.16,    2.16,    2.16,
  2.2,     2.2,     2.2,     2.2,
  2.99,    2.99,    2.99,    2.99,
  2.89,    2.89,    2.89,    2.89,
  2.94,    2.94,    2.94,    2.94,
  2.43,    2.43,    2.43,    2.43,
  2.11,    2.11,    2.11,    2.11,
  1.71,    1.71,    1.71,    1.71,
  2.25,    2.25,    2.25,    2.25,
  2.22,    2.22,    2.22,    2.22,
  2.42,    2.42,    2.42,    2.42,
  2.17,    2.17,    2.17,    2.17,
  2.21,    2.21,    2.21,    2.21,
  2.149,   2.149,   2.149,   2.149,
  2.017,   2.017,   2.017,   2.017,
  2.267,   2.267,   2.267,   2.267,
  2.58,    2.58,    2.58,    2.58,
  2.409,   2.409,   2.409,   2.409,
  2.407,   2.407,   2.407,   2.407,
  2.333,   2.333,   2.333,   2.333,
  2.409,   2.409,   2.409,   2.409,
  2.414,   2.414,   2.414,   2.414,
  2.427,   2.427,   2.427,   2.427,
  2.461,   2.461,   2.461,   2.461,
  2.454,   2.454,   2.454,   2.454,
  2.391,   2.391,   2.391,   2.391,
  2.55,    2.55,    2.55,    2.55,
  2.487,   2.487,   2.487,   2.487,
  2.4,     2.4,     2.4,     2.4,
  2.647,   2.647,   2.647,   2.647,
  2.529,   2.529,   2.529,   2.529,
  2.594,   2.594,   2.594,   2.594,
  2.477,   2.477,   2.477,   2.477,
  2.617,   2.617,   2.617,   2.617,
  2.43,    2.43,    2.43,    2.43,
  2.471,   2.471,   2.471,   2.471,
  2.604,   2.604,   2.604,   2.604,
  2.331,   2.331,   2.331,   2.331,
  2.449,   2.449,   2.449,   2.449,
  2.33,    2.33,    2.33,    2.33,
  2.39,    2.39,    2.39,    2.39,
  2.407,   2.407,   2.407,   2.407,
  2.534,   2.534,   2.534,   2.534,
  2.467,   2.467,   2.467,   2.467,
  2.414,   2.414,   2.414,   2.414,
  2.311,   2.311,   2.311,   2.311,
  2.326,   2.326,   2.326,   2.326,
  2.129,   2.129,   2.129,   2.129,
  2.029,   2.029,   2.029,   2.029,
  2.428,   2.428,   2.428,   2.428,
  2.503,   2.503,   2.503,   2.503,
  2.468,   2.468,   2.468,   2.468,
  2.596,   2.596,   2.596,   2.596,
  2.493,   2.493,   2.493,   2.493,
  2.459,   2.459,   2.459,   2.459,
  2.285,   2.285,   2.285,   2.285,
  2.257,   2.257,   2.257,   2.257,
  2.275,   2.275,   2.275,   2.275,
  2.129,   2.129,   2.129,   2.129,
  2.223,   2.223,   2.223,   2.223,
  2.186,   2.186,   2.186,   2.186,
  2.149,   2.149,   2.149,   2.149,
  2.017,   2.017,   2.017,   2.017,
  2.267,   2.267,   2.267,   2.267,
  2.58,    2.58,    2.58,    2.58,
  2.409,   2.409,   2.409,   2.409,
  2.407,   2.407,   2.407,   2.407,
  2.333,   2.333,   2.333,   2.333,
  2.409,   2.409,   2.409,   2.409,
  2.414,   2.414,   2.414,   2.414,
  2.427,   2.427,   2.427,   2.427,
  2.461,   2.461,   2.461,   2.461,
  2.454,   2.454,   2.454,   2.454,
  2.391,   2.391,   2.391,   2.391,
  2.55,    2.55,    2.55,    2.55,
  2.487,   2.487,   2.487,   2.487,
  2.4,     2.4,     2.4,     2.4,
  2.647,   2.647,   2.647,   2.647,
  2.529,   2.529,   2.529,   2.529,
  2.594,   2.594,   2.594,   2.594,
  2.477,   2.477,   2.477,   2.477,
  2.617,   2.617,   2.617,   2.617,
  2.43,    2.43,    2.43,    2.43,
  2.471,   2.471,   2.471,   2.471,
  2.604,   2.604,   2.604,   2.604,
  2.331,   2.331,   2.331,   2.331,
  2.449,   2.449,   2.449,   2.449,
  2.33,    2.33,    2.33,    2.33,
  2.39,    2.39,    2.39,    2.39,
  2.407,   2.407,   2.407,   2.407,
  2.534,   2.534,   2.534,   2.534,
  2.467,   2.467,   2.467,   2.467,
  2.414,   2.414,   2.414,   2.414,
  2.311,   2.311,   2.311,   2.311,
  2.326,   2.326,   2.326,   2.326,
  2.129,   2.129,   2.129,   2.129,
  2.029,   2.029,   2.029,   2.029,
  4.02,    4.02,    4.02,    4.02,
  3.46,    3.46,    3.46,    3.46,
  3.68,    3.68,    3.68,    3.68,
  3.94,    3.94,    3.94,    3.94,
  4.69,    4.69,    4.69,    4.69,
  4.63,    4.63,    4.63,    4.63,
  2.285,   2.285,   2.285,   2.285,
  2.257,   2.257,   2.257,   2.257,
  2.275,   2.275,   2.275,   2.275,
  2.129,   2.129,   2.129,   2.129,
  2.223,   2.223,   2.223,   2.223,
  2.186,   2.186,   2.186,   2.186,
  2.149,   2.149,   2.149,   2.149,
  2.017,   2.017,   2.017,   2.017,
  2.267,   2.267,   2.267,   2.267,
  2.58,    2.58,    2.58,    2.58,
  2.409,   2.409,   2.409,   2.409,
  2.407,   2.407,   2.407,   2.407,
  2.333,   2.333,   2.333,   2.333,
  2.409,   2.409,   2.409,   2.409,
  2.414,   2.414,   2.414,   2.414,
  2.427,   2.427,   2.427,   2.427,
  2.461,   2.461,   2.461,   2.461,
  2.454,   2.454,   2.454,   2.454,
  2.391,   2.391,   2.391,   2.391,
  2.55,    2.55,    2.55,    2.55,
  2.487,   2.487,   2.487,   2.487,
  2.4,     2.4,     2.4,     2.4,
  2.647,   2.647,   2.647,   2.647,
  2.529,   2.529,   2.529,   2.529,
  2.594,   2.594,   2.594,   2.594,
  2.477,   2.477,   2.477,   2.477,
  2.617,   2.617,   2.617,   2.617,
  2.43,    2.43,    2.43,    2.43,
  2.471,   2.471,   2.471,   2.471,
  2.604,   2.604,   2.604,   2.604,
  2.331,   2.331,   2.331,   2.331,
  2.449,   2.449,   2.449,   2.449,
  2.33,    2.33,    2.33,    2.33,
  2.39,    2.39,    2.39,    2.39,
  2.407,   2.407,   2.407,   2.407,
  2.534,   2.534,   2.534,   2.534,
  2.467,   2.467,   2.467,   2.467,
  2.414,   2.414,   2.414,   2.414,
  2.311,   2.311,   2.311,   2.311,
  2.326,   2.326,   2.326,   2.326,
  2.129,   2.129,   2.129,   2.129,
  2.029,   2.029,   2.029,   2.029,
  2.428,   2.428,   2.428,   2.428,
  2.503,   2.503,   2.503,   2.503,
  2.468,   2.468,   2.468,   2.468,
  2.596,   2.596,   2.596,   2.596,
  2.493,   2.493,   2.493,   2.493,
  2.459,   2.459,   2.459,   2.459,
  2.285,   2.285,   2.285,   2.285,
  2.257,   2.257,   2.257,   2.257,
  2.275,   2.275,   2.275,   2.275,
  2.129,   2.129,   2.129,   2.129,
  2.223,   2.223,   2.223,   2.223,
  2.186,   2.186,   2.186,   2.186,
  2.149,   2.149,   2.149,   2.149,
  2.017,   2.017,   2.017,   2.017,
  2.267,   2.267,   2.267,   2.267,
  2.58,    2.58,    2.58,    2.58,
  2.409,   2.409,   2.409,   2.409,
  2.407,   2.407,   2.407,   2.407,
  2.333,   2.333,   2.333,   2.333,
  2.409,   2.409,   2.409,   2.409,
  2.414,   2.414,   2.414,   2.414,
  2.427,   2.427,   2.427,   2.427,
  2.461,   2.461,   2.461,   2.461,
  2.454,   2.454,   2.454,   2.454,
  2.391,   2.391,   2.391,   2.391,
  2.55,    2.55,    2.55,    2.55,
  2.487,   2.487,   2.487,   2.487,
  2.4,     2.4,     2.4,     2.4,
  2.647,   2.647,   2.647,   2.647,
  2.529,   2.529,   2.529,   2.529,
  2.594,   2.594,   2.594,   2.594,
  2.477,   2.477,   2.477,   2.477,
  2.617,   2.617,   2.617,   2.617,
  2.43,    2.43,    2.43,    2.43,
  2.471,   2.471,   2.471,   2.471,
  2.604,   2.604,   2.604,   2.604,
  2.331,   2.331,   2.331,   2.331,
  2.449,   2.449,   2.449,   2.449,
  2.33,    2.33,    2.33,    2.33,
  2.39,    2.39,    2.39,    2.39,
  2.407,   2.407,   2.407,   2.407,
  2.534,   2.534,   2.534,   2.534,
  2.467,   2.467,   2.467,   2.467,
  2.414,   2.414,   2.414,   2.414,
  2.311,   2.311,   2.311,   2.311,
  2.326,   2.326,   2.326,   2.326,
  2.129,   2.129,   2.129,   2.129,
  2.029,   2.029,   2.029,   2.029,
  2.428,   2.428,   2.428,   2.428,
  2.503,   2.503,   2.503,   2.503,
  2.468,   2.468,   2.468,   2.468,
  2.596,   2.596,   2.596,   2.596,
  2.493,   2.493,   2.493,   2.493,
  2.459,   2.459,   2.459,   2.459,
  2.285,   2.285,   2.285,   2.285,
  2.257,   2.257,   2.257,   2.257,
  2.275,   2.275,   2.275,   2.275,
  2.129,   2.129,   2.129,   2.129,
  2.223,   2.223,   2.223,   2.223,
  2.186,   2.186,   2.186,   2.186,
  2.149,   2.149,   2.149,   2.149,
  2.017,   2.017,   2.017,   2.017,
  2.267,   2.267,   2.267,   2.267,
  2.58,    2.58,    2.58,    2.58,
  2.409,   2.409,   2.409,   2.409,
  2.407,   2.407,   2.407,   2.407,
  2.333,   2.333,   2.333,   2.333,
  2.409,   2.409,   2.409,   2.409,
  2.414,   2.414,   2.414,   2.414,
  2.427,   2.427,   2.427,   2.427,
  2.461,   2.461,   2.461,   2.461,
  2.454,   2.454,   2.454,   2.454,
  2.391,   2.391,   2.391,   2.391,
  2.55,    2.55,    2.55,    2.55,
  2.487,   2.487,   2.487,   2.487,
  2.4,     2.4,     2.4,     2.4,
  2.647,   2.647,   2.647,   2.647,
  2.529,   2.529,   2.529,   2.529,
  2.594,   2.594,   2.594,   2.594,
  2.477,   2.477,   2.477,   2.477,
  2.617,   2.617,   2.617,   2.617,
  2.43,    2.43,    2.43,    2.43,
  2.471,   2.471,   2.471,   2.471,
  2.604,   2.604,   2.604,   2.604,
  2.331,   2.331,   2.331,   2.331,
  2.449,   2.449,   2.449,   2.449,
  2.33,    2.33,    2.33,    2.33,
  2.39,    2.39,    2.39,    2.39,
  2.407,   2.407,   2.407,   2.407,
  2.534,   2.534,   2.534,   2.534,
  2.467,   2.467,   2.467,   2.467,
  2.414,   2.414,   2.414,   2.414,
  2.311,   2.311,   2.311,   2.311,
  2.326,   2.326,   2.326,   2.326,
  2.129,   2.129,   2.129,   2.129,
  2.029,   2.029,   2.029,   2.029,
  2.428,   2.428,   2.428,   2.428,
  2.503,   2.503,   2.503,   2.503,
  2.468,   2.468,   2.468,   2.468,
  2.596,   2.596,   2.596,   2.596,
  2.493,   2.493,   2.493,   2.493,
  2.459,   2.459,   2.459,   2.459,
  2.285,   2.285,   2.285,   2.285,
  2.257,   2.257,   2.257,   2.257,
  2.275,   2.275,   2.275,   2.275,
  2.129,   2.129,   2.129,   2.129,
  2.223,   2.223,   2.223,   2.223,
  2.186,   2.186,   2.186,   2.186,
  2.149,   2.149,   2.149,   2.149,
  2.017,   2.017,   2.017,   2.017,
  2.267,   2.267,   2.267,   2.267,
  2.58,    2.58,    2.58,    2.58,
  2.409,   2.409,   2.409,   2.409,
  2.407,   2.407,   2.407,   2.407,
  2.333,   2.333,   2.333,   2.333,
  2.409,   2.409,   2.409,   2.409,
  2.414,   2.414,   2.414,   2.414,
  2.427,   2.427,   2.427,   2.427,
  2.461,   2.461,   2.461,   2.461,
  2.454,   2.454,   2.454,   2.454,
  2.391,   2.391,   2.391,   2.391,
  2.55,    2.55,    2.55,    2.55,
  2.487,   2.487,   2.487,   2.487,
  2.4,     2.4,     2.4,     2.4,
  2.647,   2.647,   2.647,   2.647,
  2.529,   2.529,   2.529,   2.529,
  2.594,   2.594,   2.594,   2.594,
  2.477,   2.477,   2.477,   2.477,
  2.617,   2.617,   2.617,   2.617,
  2.43,    2.43,    2.43,    2.43,
  2.471,   2.471,   2.471,   2.471,
  2.604,   2.604,   2.604,   2.604,
  2.331,   2.331,   2.331,   2.331,
  2.449,   2.449,   2.449,   2.449,
  2.33,    2.33,    2.33,    2.33,
  2.39,    2.39,    2.39,    2.39,
  2.407,   2.407,   2.407,   2.407,
  2.534,   2.534,   2.534,   2.534,
  2.467,   2.467,   2.467,   2.467,
  2.414,   2.414,   2.414,   2.414,
  2.311,   2.311,   2.311,   2.311,
  2.326,   2.326,   2.326,   2.326,
  2.129,   2.129,   2.129,   2.129,
  2.029,   2.029,   2.029,   2.029,
  2.428,   2.428,   2.428,   2.428,
  2.503,   2.503,   2.503,   2.503,
  2.468,   2.468,   2.468,   2.468,
  2.596,   2.596,   2.596,   2.596,
  2.493,   2.493,   2.493,   2.493,
  2.459,   2.459,   2.459,   2.459,
  2.285,   2.285,   2.285,   2.285,
  2.257,   2.257,   2.257,   2.257,
  2.275,   2.275,   2.275,   2.275,
  2.129,   2.129,   2.129,   2.129,
  2.223,   2.223,   2.223,   2.223,
  2.186,   2.186,   2.186,   2.186,
  2.149,   2.149,   2.149,   2.149,
  2.017,   2.017,   2.017,   2.017,
  2.267,   2.267,   2.267,   2.267,
  2.58,    2.58,    2.58,    2.58,
  2.409,   2.409,   2.409,   2.409,
  2.407,   2.407,   2.407,   2.407,
  2.333,   2.333,   2.333,   2.333,
  2.409,   2.409,   2.409,   2.409,
  2.414,   2.414,   2.414,   2.414,
  2.427,   2.427,   2.427,   2.427,
  2.461,   2.461,   2.461,   2.461,
  2.454,   2.454,   2.454,   2.454,
  2.391,   2.391,   2.391,   2.391,
  2.55,    2.55,    2.55,    2.55,
  2.487,   2.487,   2.487,   2.487,
  2.4,     2.4,     2.4,     2.4,
  2.647,   2.647,   2.647,   2.647,
  2.529,   2.529,   2.529,   2.529,
  2.594,   2.594,   2.594,   2.594,
  2.477,   2.477,   2.477,   2.477,
  2.617,   2.617,   2.617,   2.617,
  2.43,    2.43,    2.43,    2.43,
  2.471,   2.471,   2.471,   2.471,
  2.604,   2.604,   2.604,   2.604,
  2.331,   2.331,   2.331,   2.331,
  2.449,   2.449,   2.449,   2.449,
  2.33,    2.33,    2.33,    2.33,
  2.39,    2.39,    2.39,    2.39,
  2.407,   2.407,   2.407,   2.407,
  2.534,   2.534,   2.534,   2.534,
  2.467,   2.467,   2.467,   2.467,
  2.414,   2.414,   2.414,   2.414,
  2.311,   2.311,   2.311,   2.311,
  3.1,     3.1,     3.1,     3.1,
  2.34,    2.34,    2.34,    2.34,
  2.27,    2.27,    2.27,    2.27,
  2.84,    2.84,    2.84,    2.84,
  2.72,    2.72,    2.72,    2.72,
  2.32,    2.32,    2.32,    2.32,
  2.21,    2.21,    2.21,    2.21,
  2.26,    2.26,    2.26,    2.26,
  2.17,    2.17,    2.17,    2.17,
  2.86,    2.86,    2.86,    2.86,
  2.73,    2.73,    2.73,    2.73,
  2.61,    2.61,    2.61,    2.61,
  2.04,    2.04,    2.04,    2.04,
  1.32,    1.32,    1.32,    1.32,
  1.75,    1.75,    1.75,    1.75,
  2.14,    2.14,    2.14,    2.14,
  2.26,    2.26,    2.26,    2.26,
  2.32,    2.32,    2.32,    2.32,
  3.1,     3.1,     3.1,     3.1,
  2.47,    2.47,    2.47,    2.47,
  3.07,    3.07,    3.07,    3.07,
  2.96,    2.96,    2.96,    2.96,
  2.29,    2.29,    2.29,    2.29,
  1.89,    1.89,    1.89,    1.89,
  1.61,    1.61,    1.61,    1.61,
  1.9,     1.9,     1.9,     1.9,
  1.94,    1.94,    1.94,    1.94,
  1.25,    1.25,    1.25,    1.25,
  1.5,     1.5,     1.5,     1.5,
  2.34,    2.34,    2.34,    2.34,
  2.25,    2.25,    2.25,    2.25,
  2.7,     2.7,     2.7,     2.7,
  2.81,    2.81,    2.81,    2.81,
  2.97,    2.97,    2.97,    2.97,
  2.54,    2.54,    2.54,    2.54,
  2.97,    2.97,    2.97,    2.97,
  2.88,    2.88,    2.88,    2.88,
  2.25,    2.25,    2.25,    2.25,
  3.41,    3.41,    3.41,    3.41,
  2.64,    2.64,    2.64,    2.64,
  2.48,    2.48,    2.48,    2.48,
  2.41,    2.41,    2.41,    2.41,
  2.65,    2.65,    2.65,    2.65,
  2.76,    2.76,    2.76,    2.76,
  3.04,    3.04,    3.04,    3.04,
  3.33,    3.33,    3.33,    3.33,
  3.04,    3.04,    3.04,    3.04,
  2.69,    2.69,    2.69,    2.69,
  2.74,    2.74,    2.74,    2.74,
  2.69,    2.69,    2.69,    2.69,
  2.19,    2.19,    2.19,    2.19,
  2.38,    2.38,    2.38,    2.38,
  2.6,     2.6,     2.6,     2.6,
  3.05,    3.05,    3.05,    3.05,
  3.85,    3.85,    3.85,    3.85,
  2.97,    2.97,    2.97,    2.97,
  2.97,    2.97,    2.97,    2.97,
  3.31,    3.31,    3.31,    3.31,
  2.71,    2.71,    2.71,    2.71,
  2.84,    2.84,    2.84,    2.84,
  2.76,    2.76,    2.76,    2.76,
  3.39,    3.39,    3.39,    3.39,
  2.74,    2.74,    2.74,    2.74,
  2.37,    2.37,    2.37,    2.37,
  2.04,    2.04,    2.04,    2.04,
  2.22,    2.22,    2.22,    2.22,
  2.9,     2.9,     2.9,     2.9,
  2.06,    2.06,    2.06,    2.06,
  2.56,    2.56,    2.56,    2.56,
  2.39,    2.39,    2.39,    2.39,
  2.89,    2.89,    2.89,    2.89,
  2.4,     2.4,     2.4,     2.4,
  2.63,    2.63,    2.63,    2.63,
  3.14,    3.14,    3.14,    3.14,
  2.66,    2.66,    2.66,    2.66,
  2.89,    2.89,    2.89,    2.89,
  2.78,    2.78,    2.78,    2.78,
  2.17,    2.17,    2.17,    2.17,
  2.46,    2.46,    2.46,    2.46,
  2.73,    2.73,    2.73,    2.73,
  2.7,     2.7,     2.7,     2.7,
  2.93,    2.93,    2.93,    2.93,
  2.61,    2.61,    2.61,    2.61,
  2.26,    2.26,    2.26,    2.26,
  2.43,    2.43,    2.43,    2.43,
  2.25,    2.25,    2.25,    2.25,
  2,       2,       2,       2,
  1.14,    1.14,    1.14,    1.14,
  1.56,    1.56,    1.56,    1.56,
  1.27,    1.27,    1.27,    1.27,
  1.7,     1.7,     1.7,     1.7,
  1.8,     1.8,     1.8,     1.8,
  1.43,    1.43,    1.43,    1.43,
  1.22,    1.22,    1.22,    1.22,
  1.41,    1.41,    1.41,    1.41,
  1.46,    1.46,    1.46,    1.46,
  1.04,    1.04,    1.04,    1.04,
  0.97,    0.97,    0.97,    0.97,
  1.04,    1.04,    1.04,    1.04,
  0.77,    0.77,    0.77,    0.77,
  1.06,    1.06,    1.06,    1.06,
  0.83,    0.83,    0.83,    0.83,
  1.25,    1.25,    1.25,    1.25,
  1.21,    1.21,    1.21,    1.21,
  0.74,    0.74,    0.74,    0.74,
  1.1,     1.1,     1.1,     1.1,
  0.99,    0.99,    0.99,    0.99,
  1.29,    1.29,    1.29,    1.29,
  1.08,    1.08,    1.08,    1.08,
  1.27,    1.27,    1.27,    1.27,
  1.09,    1.09,    1.09,    1.09,
  0.79,    0.79,    0.79,    0.79,
  0.76,    0.76,    0.76,    0.76,
  0.87,    0.87,    0.87,    0.87,
  1,       1,       1,       1,
  1.19,    1.19,    1.19,    1.19,
  0.99,    0.99,    0.99,    0.99,
  1.06,    1.06,    1.06,    1.06,
  1.08,    1.08,    1.08,    1.08,
  1.23,    1.23,    1.23,    1.23,
  1.09,    1.09,    1.09,    1.09,
  1.19,    1.19,    1.19,    1.19,
  1.56,    1.56,    1.56,    1.56,
  1.43,    1.43,    1.43,    1.43,
  1.68,    1.68,    1.68,    1.68,
  1.77,    1.77,    1.77,    1.77,
  1.74,    1.74,    1.74,    1.74,
  1.76,    1.76,    1.76,    1.76,
  1.44,    1.44,    1.44,    1.44,
  1.45,    1.45,    1.45,    1.45,
  1.46,    1.46,    1.46,    1.46,
  1.55,    1.55,    1.55,    1.55,
  1.56,    1.56,    1.56,    1.56,
  1.59,    1.59,    1.59,    1.59,
  1.74,    1.74,    1.74,    1.74,
  1.59,    1.59,    1.59,    1.59,
  2.06,    2.06,    2.06,    2.06,
  1.79,    1.79,    1.79,    1.79,
  1.7,     1.7,     1.7,     1.7,
  1.57,    1.57,    1.57,    1.57,
  1.94,    1.94,    1.94,    1.94,
  2.2,     2.2,     2.2,     2.2,
  1.85,    1.85,    1.85,    1.85,
  2.13,    2.13,    2.13,    2.13,
  2.2,     2.2,     2.2,     2.2,
  1.8,     1.8,     1.8,     1.8,
  1.93,    1.93,    1.93,    1.93,
  2.45,    2.45,    2.45,    2.45,
  2.27,    2.27,    2.27,    2.27,
  2.18,    2.18,    2.18,    2.18,
  2.21,    2.21,    2.21,    2.21,
  1.56,    1.56,    1.56,    1.56,
  1.78,    1.78,    1.78,    1.78,
  1.86,    1.86,    1.86,    1.86,
  1.76,    1.76,    1.76,    1.76,
  1.98,    1.98,    1.98,    1.98,
  2.09,    2.09,    2.09,    2.09,
  2.51,    2.51,    2.51,    2.51,
  2.42,    2.42,    2.42,    2.42,
  2.37,    2.37,    2.37,    2.37,
  2.27,    2.27,    2.27,    2.27,
  2.26,    2.26,    2.26,    2.26,
  2.28,    2.28,    2.28,    2.28,
  2.37,    2.37,    2.37,    2.37,
  2.08,    2.08,    2.08,    2.08,
  2.05,    2.05,    2.05,    2.05,
  2.55,    2.55,    2.55,    2.55,
  2.55,    2.55,    2.55,    2.55,
  2.69,    2.69,    2.69,    2.69,
  2.52,    2.52,    2.52,    2.52,
  2.96,    2.96,    2.96,    2.96,
  3.21,    3.21,    3.21,    3.21,
  3.03,    3.03,    3.03,    3.03,
  2.57,    2.57,    2.57,    2.57,
  2.44,    2.44,    2.44,    2.44,
  2.73,    2.73,    2.73,    2.73,
  2.87,    2.87,    2.87,    2.87,
  2.83,    2.83,    2.83,    2.83,
  3,       3,       3,       3,
  2.98,    2.98,    2.98,    2.98,
  2.57,    2.57,    2.57,    2.57,
  2.66,    2.66,    2.66,    2.66,
  2.95,    2.95,    2.95,    2.95,
  2.81,    2.81,    2.81,    2.81,
  2.76,    2.76,    2.76,    2.76,
  2.49,    2.49,    2.49,    2.49,
  3.03,    3.03,    3.03,    3.03,
  2.83,    2.83,    2.83,    2.83,
  2.9,     2.9,     2.9,     2.9,
  2.61,    2.61,    2.61,    2.61,
  3.01,    3.01,    3.01,    3.01,
  2.56,    2.56,    2.56,    2.56,
  2.47,    2.47,    2.47,    2.47,
  3.04,    3.04,    3.04,    3.04,
  2.46,    2.46,    2.46,    2.46,
  2.63,    2.63,    2.63,    2.63,
  2.67,    2.67,    2.67,    2.67,
  2.74,    2.74,    2.74,    2.74,
  2.56,    2.56,    2.56,    2.56,
  2.55,    2.55,    2.55,    2.55,
  3.06,    3.06,    3.06,    3.06,
  2.98,    2.98,    2.98,    2.98,
  2.77,    2.77,    2.77,    2.77,
  2.59,    2.59,    2.59,    2.59,
  2.25,    2.25,    2.25,    2.25,
  2.48,    2.48,    2.48,    2.48,
  2.53,    2.53,    2.53,    2.53,
  2.68,    2.68,    2.68,    2.68,
  2.65,    2.65,    2.65,    2.65,
  2.58,    2.58,    2.58,    2.58,
  2.47,    2.47,    2.47,    2.47,
  2.13,    2.13,    2.13,    2.13,
  2.26,    2.26,    2.26,    2.26,
  2.14,    2.14,    2.14,    2.14,
  1.96,    1.96,    1.96,    1.96,
  2.31,    2.31,    2.31,    2.31,
  2.39,    2.39,    2.39,    2.39,
  2.25,    2.25,    2.25,    2.25,
  1.89,    1.89,    1.89,    1.89,
  1.98,    1.98,    1.98,    1.98,
  2.31,    2.31,    2.31,    2.31,
  2.14,    2.14,    2.14,    2.14,
  2.07,    2.07,    2.07,    2.07,
  2.51,    2.51,    2.51,    2.51,
  2.24,    2.24,    2.24,    2.24,
  2.45,    2.45,    2.45,    2.45,
  2.67,    2.67,    2.67,    2.67,
  3.04,    3.04,    3.04,    3.04,
  2.58,    2.58,    2.58,    2.58,
  2.77,    2.77,    2.77,    2.77,
  2.88,    2.88,    2.88,    2.88,
  3.21,    3.21,    3.21,    3.21,
  3.79,    3.79,    3.79,    3.79,
  3.11,    3.11,    3.11,    3.11,
  2.59,    2.59,    2.59,    2.59,
  2.95,    2.95,    2.95,    2.95,
  2.63,    2.63,    2.63,    2.63,
  2.42,    2.42,    2.42,    2.42,
  2.42,    2.42,    2.42,    2.42,
  2.38,    2.38,    2.38,    2.38,
  2.24,    2.24,    2.24,    2.24,
  2.22,    2.22,    2.22,    2.22,
  2.07,    2.07,    2.07,    2.07,
  2.11,    2.11,    2.11,    2.11,
  2.17,    2.17,    2.17,    2.17,
  2.09,    2.09,    2.09,    2.09,
  2.22,    2.22,    2.22,    2.22,
  2.41,    2.41,    2.41,    2.41,
  2.28,    2.28,    2.28,    2.28,
  2.15,    2.15,    2.15,    2.15,
  2.18,    2.18,    2.18,    2.18,
  2.11,    2.11,    2.11,    2.11,
  2.23,    2.23,    2.23,    2.23,
  2.32,    2.32,    2.32,    2.32,
  2.27,    2.27,    2.27,    2.27,
  2.05,    2.05,    2.05,    2.05,
  2.12,    2.12,    2.12,    2.12,
  1.85,    1.85,    1.85,    1.85,
  2.02,    2.02,    2.02,    2.02,
  2.22,    2.22,    2.22,    2.22,
  1.81,    1.81,    1.81,    1.81,
  2,       2,       2,       2,
  2.09,    2.09,    2.09,    2.09,
  2.16,    2.16,    2.16,    2.16,
  2.2,     2.2,     2.2,     2.2,
  2.31,    2.31,    2.31,    2.31,
  2.01,    2.01,    2.01,    2.01,
  1.91,    1.91,    1.91,    1.91,
  2.08,    2.08,    2.08,    2.08,
  2.22,    2.22,    2.22,    2.22,
  1.89,    1.89,    1.89,    1.89,
  2.11,    2.11,    2.11,    2.11,
  1.9,     1.9,     1.9,     1.9,
  1.92,    1.92,    1.92,    1.92,
  2.05,    2.05,    2.05,    2.05,
  2.38,    2.38,    2.38,    2.38,
  2.1,     2.1,     2.1,     2.1,
  2.18,    2.18,    2.18,    2.18,
  2.01,    2.01,    2.01,    2.01,
  1.79,    1.79,    1.79,    1.79,
  1.2,     1.2,     1.2,     1.2,
  1.24,    1.24,    1.24,    1.24,
  1.97,    1.97,    1.97,    1.97,
  1.86,    1.86,    1.86,    1.86,
  1.94,    1.94,    1.94,    1.94,
  2,       2,       2,       2,
  1.81,    1.81,    1.81,    1.81,
  1.77,    1.77,    1.77,    1.77,
  1.66,    1.66,    1.66,    1.66,
  1.82,    1.82,    1.82,    1.82,
  2.11,    2.11,    2.11,    2.11,
  2.45,    2.45,    2.45,    2.45,
  2.59,    2.59,    2.59,    2.59,
  2.43,    2.43,    2.43,    2.43,
  2.18,    2.18,    2.18,    2.18,
  2.36,    2.36,    2.36,    2.36,
  2.39,    2.39,    2.39,    2.39,
  2.31,    2.31,    2.31,    2.31,
  2.67,    2.67,    2.67,    2.67,
  2.56,    2.56,    2.56,    2.56,
  2.16,    2.16,    2.16,    2.16,
  2.32,    2.32,    2.32,    2.32,
  2.48,    2.48,    2.48,    2.48,
  2.64,    2.64,    2.64,    2.64,
  2.88,    2.88,    2.88,    2.88,
  2.28,    2.28,    2.28,    2.28,
  2.16,    2.16,    2.16,    2.16,
  2.12,    2.12,    2.12,    2.12,
  2.27,    2.27,    2.27,    2.27,
  2.22,    2.22,    2.22,    2.22,
  2.5,     2.5,     2.5,     2.5,
  2.35,    2.35,    2.35,    2.35,
  2.49,    2.49,    2.49,    2.49,
  2.09,    2.09,    2.09,    2.09,
  2.27,    2.27,    2.27,    2.27,
  2.25,    2.25,    2.25,    2.25,
  2.28,    2.28,    2.28,    2.28,
  2.07,    2.07,    2.07,    2.07,
  2.49,    2.49,    2.49,    2.49,
  2.44,    2.44,    2.44,    2.44,
  2.16,    2.16,    2.16,    2.16,
  2.33,    2.33,    2.33,    2.33,
  1.67,    1.67,    1.67,    1.67,
  1.75,    1.75,    1.75,    1.75,
  1.75,    1.75,    1.75,    1.75,
  1.873,   1.873,   1.873,   1.873,
  1.21,    1.21,    1.21,    1.21,
  1.81,    1.81,    1.81,    1.81,
  2.3,     2.3,     2.3,     2.3,
  2.02,    2.02,    2.02,    2.02,
  2.53,    2.53,    2.53,    2.53,
  1.63,    1.63,    1.63,    1.63,
  1.31,    1.31,    1.31,    1.31,
  1.65,    1.65,    1.65,    1.65,
  1.35,    1.35,    1.35,    1.35,
  1.19,    1.19,    1.19,    1.19,
  1.35,    1.35,    1.35,    1.35,
  1.83,    1.83,    1.83,    1.83,
  1.87,    1.87,    1.87,    1.87,
  2.25,    2.25,    2.25,    2.25,
  2.59,    2.59,    2.59,    2.59,
  2.38,    2.38,    2.38,    2.38,
  2.34,    2.34,    2.34,    2.34,
  1.92,    1.92,    1.92,    1.92,
  1.62,    1.62,    1.62,    1.62,
  2.11,    2.11,    2.11,    2.11,
  2.74,    2.74,    2.74,    2.74,
  2.52,    2.52,    2.52,    2.52,
  2.08,    2.08,    2.08,    2.08,
  2.04,    2.04,    2.04,    2.04,
  1.97,    1.97,    1.97,    1.97,
  2.06,    2.06,    2.06,    2.06,
  2.27,    2.27,    2.27,    2.27,
  2.08,    2.08,    2.08,    2.08,
  2.05,    2.05,    2.05,    2.05,
  1.79,    1.79,    1.79,    1.79,
  1.94,    1.94,    1.94,    1.94,
  2.19,    2.19,    2.19,    2.19,
  2.18,    2.18,    2.18,    2.18,
  2.37,    2.37,    2.37,    2.37,
  2.53,    2.53,    2.53,    2.53,
  2.36,    2.36,    2.36,    2.36,
  2.3,     2.3,     2.3,     2.3,
  2.33,    2.33,    2.33,    2.33,
  2.22,    2.22,    2.22,    2.22,
  2.33,    2.33,    2.33,    2.33,
  2.16,    2.16,    2.16,    2.16,
  2.24,    2.24,    2.24,    2.24,
  2.13,    2.13,    2.13,    2.13,
  2.2,     2.2,     2.2,     2.2,
  1.97,    1.97,    1.97,    1.97,
  1.76,    1.76,    1.76,    1.76,
  1.79,    1.79,    1.79,    1.79,
  1.7,     1.7,     1.7,     1.7,
  1.32,    1.32,    1.32,    1.32,
  1.46,    1.46,    1.46,    1.46,
  1.24,    1.24,    1.24,    1.24,
  1.38,    1.38,    1.38,    1.38,
  0.97,    0.97,    0.97,    0.97,
  1.39,    1.39,    1.39,    1.39,
  1.07,    1.07,    1.07,    1.07,
  1.1,     1.1,     1.1,     1.1,
  1.5,     1.5,     1.5,     1.5,
  1.28,    1.28,    1.28,    1.28,
  1.63,    1.63,    1.63,    1.63,
  1.86,    1.86,    1.86,    1.86,
  2.26,    2.26,    2.26,    2.26,
  2.37,    2.37,    2.37,    2.37,
  2.46,    2.46,    2.46,    2.46,
  2.25,    2.25,    2.25,    2.25,
  2.17,    2.17,    2.17,    2.17,
  2.23,    2.23,    2.23,    2.23,
  2.12,    2.12,    2.12,    2.12,
  2.56,    2.56,    2.56,    2.56,
  2.56,    2.56,    2.56,    2.56,
  2.22,    2.22,    2.22,    2.22,
  2.24,    2.24,    2.24,    2.24,
  2.83,    2.83,    2.83,    2.83,
  2.76,    2.76,    2.76,    2.76,
  2.86,    2.86,    2.86,    2.86,
  2.49,    2.49,    2.49,    2.49,
  2.74,    2.74,    2.74,    2.74,
  2.49,    2.49,    2.49,    2.49,
  2.31,    2.31,    2.31,    2.31,
  2.76,    2.76,    2.76,    2.76,
  2.38,    2.38,    2.38,    2.38,
  2.34,    2.34,    2.34,    2.34,
  2.57,    2.57,    2.57,    2.57,
  2.26,    2.26,    2.26,    2.26,
  2.42,    2.42,    2.42,    2.42,
  2.4,     2.4,     2.4,     2.4,
  2.42,    2.42,    2.42,    2.42,
  2.68,    2.68,    2.68,    2.68,
  2.88,    2.88,    2.88,    2.88,
  2.67,    2.67,    2.67,    2.67,
  2.3,     2.3,     2.3,     2.3,
  2.31,    2.31,    2.31,    2.31,
  2.21,    2.21,    2.21,    2.21,
  2.88,    2.88,    2.88,    2.88,
  2.73,    2.73,    2.73,    2.73,
  2.24,    2.24,    2.24,    2.24,
  2.28,    2.28,    2.28,    2.28,
  2.31,    2.31,    2.31,    2.31,
  2.69,    2.69,    2.69,    2.69,
  3.21,    3.21,    3.21,    3.21,
  3.09,    3.09,    3.09,    3.09,
  2.89,    2.89,    2.89,    2.89,
  2.76,    2.76,    2.76,    2.76,
  3.64,    3.64,    3.64,    3.64,
  3.37,    3.37,    3.37,    3.37,
  2.79,    2.79,    2.79,    2.79,
  2.73,    2.73,    2.73,    2.73,
  2.63,    2.63,    2.63,    2.63,
  2.82,    2.82,    2.82,    2.82,
  2.56,    2.56,    2.56,    2.56,
  2.79,    2.79,    2.79,    2.79,
  3.12,    3.12,    3.12,    3.12,
  3.13,    3.13,    3.13,    3.13,
  2.99,    2.99,    2.99,    2.99,
  3.27,    3.27,    3.27,    3.27,
  3.03,    3.03,    3.03,    3.03,
  3.08,    3.08,    3.08,    3.08,
  2.5,     2.5,     2.5,     2.5,
  2.95,    2.95,    2.95,    2.95,
  2.84,    2.84,    2.84,    2.84,
  2.99,    2.99,    2.99,    2.99,
  2.87,    2.87,    2.87,    2.87,
  2.46,    2.46,    2.46,    2.46,
  2.88,    2.88,    2.88,    2.88,
  2.4,     2.4,     2.4,     2.4,
  3.22,    3.22,    3.22,    3.22,
  3.1,     3.1,     3.1,     3.1,
  2.89,    2.89,    2.89,    2.89,
  3.28,    3.28,    3.28,    3.28,
  3.24,    3.24,    3.24,    3.24,
  2.74,    2.74,    2.74,    2.74,
  2.77,    2.77,    2.77,    2.77,
  2.5,     2.5,     2.5,     2.5,
  2.22,    2.22,    2.22,    2.22,
  2.18,    2.18,    2.18,    2.18,
  2.28,    2.28,    2.28,    2.28,
  2.18,    2.18,    2.18,    2.18,
  1.59,    1.59,    1.59,    1.59,
  1.79,    1.79,    1.79,    1.79,
  1.85,    1.85,    1.85,    1.85,
  1.99,    1.99,    1.99,    1.99,
  1.9,     1.9,     1.9,     1.9,
  2.27,    2.27,    2.27,    2.27,
  2.26,    2.26,    2.26,    2.26,
  2.37,    2.37,    2.37,    2.37,
  2.53,    2.53,    2.53,    2.53,
  2.39,    2.39,    2.39,    2.39,
  2.4,     2.4,     2.4,     2.4,
  2.29,    2.29,    2.29,    2.29,
  2.14,    2.14,    2.14,    2.14,
  1.65,    1.65,    1.65,    1.65,
  1.98,    1.98,    1.98,    1.98,
  1.71,    1.71,    1.71,    1.71,
  1.59,    1.59,    1.59,    1.59,
  1.73,    1.73,    1.73,    1.73,
  1.59,    1.59,    1.59,    1.59,
  1.48,    1.48,    1.48,    1.48,
  1.33,    1.33,    1.33,    1.33,
  1.24,    1.24,    1.24,    1.24,
  1.39,    1.39,    1.39,    1.39,
  1.57,    1.57,    1.57,    1.57,
  1.56,    1.56,    1.56,    1.56,
  1.71,    1.71,    1.71,    1.71,
  1.49,    1.49,    1.49,    1.49,
  1.63,    1.63,    1.63,    1.63,
  1.29,    1.29,    1.29,    1.29,
  1,       1,       1,       1,
  1.38,    1.38,    1.38,    1.38,
  1.43,    1.43,    1.43,    1.43,
  1.42,    1.42,    1.42,    1.42,
  1.76,    1.76,    1.76,    1.76,
  2.78,    2.78,    2.78,    2.78,
  2.58,    2.58,    2.58,    2.58,
  3.01,    3.01,    3.01,    3.01,
  2.69,    2.69,    2.69,    2.69,
  3.02,    3.02,    3.02,    3.02,
  2.98,    2.98,    2.98,    2.98,
  3.18,    3.18,    3.18,    3.18,
  2.99,    2.99,    2.99,    2.99,
  2.94,    2.94,    2.94,    2.94,
  3.32,    3.32,    3.32,    3.32,
  3.2,     3.2,     3.2,     3.2,
  2.84,    2.84,    2.84,    2.84,
  2.61,    2.61,    2.61,    2.61,
  2.96,    2.96,    2.96,    2.96,
  3.09,    3.09,    3.09,    3.09,
  2.81,    2.81,    2.81,    2.81,
  2.4,     2.4,     2.4,     2.4,
  2.74,    2.74,    2.74,    2.74,
  2.92,    2.92,    2.92,    2.92,
  2.96,    2.96,    2.96,    2.96,
  2.78,    2.78,    2.78,    2.78,
  2.77,    2.77,    2.77,    2.77,
  2.5,     2.5,     2.5,     2.5,
  2.01,    2.01,    2.01,    2.01,
  2.37,    2.37,    2.37,    2.37,
  1.95,    1.95,    1.95,    1.95,
  1.82,    1.82,    1.82,    1.82,
  1.81,    1.81,    1.81,    1.81,
  1.68,    1.68,    1.68,    1.68,
  1.53,    1.53,    1.53,    1.53,
  1.48,    1.48,    1.48,    1.48,
  1.38,    1.38,    1.38,    1.38,
  1.46,    1.46,    1.46,    1.46,
  1.19,    1.19,    1.19,    1.19,
  1.5,     1.5,     1.5,     1.5,
  1.21,    1.21,    1.21,    1.21,
  1.34,    1.34,    1.34,    1.34,
  1.2,     1.2,     1.2,     1.2,
  1.24,    1.24,    1.24,    1.24,
  1.28,    1.28,    1.28,    1.28,
  1.13,    1.13,    1.13,    1.13,
  0.71,    0.71,    0.71,    0.71,
  0.62,    0.62,    0.62,    0.62,
  0.75,    0.75,    0.75,    0.75,
  0.61,    0.61,    0.61,    0.61,
  0.89,    0.89,    0.89,    0.89,
  0.9,     0.9,     0.9,     0.9,
  0.7,     0.7,     0.7,     0.7,
  1.17,    1.17,    1.17,    1.17,
  0.9,     0.9,     0.9,     0.9,
  0.99,    0.99,    0.99,    0.99,
  0.9,     0.9,     0.9,     0.9,
  0.85,    0.85,    0.85,    0.85,
  1.41,    1.41,    1.41,    1.41,
  1.93,    1.93,    1.93,    1.93,
  1.77,    1.77,    1.77,    1.77,
  1.37,    1.37,    1.37,    1.37,
  1.33,    1.33,    1.33,    1.33,
  1.75,    1.75,    1.75,    1.75,
  2.28,    2.28,    2.28,    2.28,
  2.21,    2.21,    2.21,    2.21,
  2.18,    2.18,    2.18,    2.18,
  1.46,    1.46,    1.46,    1.46,
  1.87,    1.87,    1.87,    1.87,
  1.79,    1.79,    1.79,    1.79,
  1.89,    1.89,    1.89,    1.89,
  1.67,    1.67,    1.67,    1.67,
  1.66,    1.66,    1.66,    1.66,
  1.71,    1.71,    1.71,    1.71,
  1.37,    1.37,    1.37,    1.37,
  1.39,    1.39,    1.39,    1.39,
  1.16,    1.16,    1.16,    1.16,
  0.9,     0.9,     0.9,     0.9,
  1.08,    1.08,    1.08,    1.08,
  0.59,    0.59,    0.59,    0.59,
  0.31,    0.31,    0.31,    0.31,
  0.67,    0.67,    0.67,    0.67,
  1.1,     1.1,     1.1,     1.1,
  0.77,    0.77,    0.77,    0.77,
  1.64,    1.64,    1.64,    1.64,
  1.04,    1.04,    1.04,    1.04,
  1.11,    1.11,    1.11,    1.11,
  0.98,    0.98,    0.98,    0.98,
  1.24,    1.24,    1.24,    1.24,
  1.31,    1.31,    1.31,    1.31,
  0.81,    0.81,    0.81,    0.81,
  0.62,    0.62,    0.62,    0.62,
  0.65,    0.65,    0.65,    0.65,
  0.76,    0.76,    0.76,    0.76,
  1.1,     1.1,     1.1,     1.1,
  1.14,    1.14,    1.14,    1.14,
  1.54,    1.54,    1.54,    1.54,
  1.2,     1.2,     1.2,     1.2,
  1.51,    1.51,    1.51,    1.51,
  1.53,    1.53,    1.53,    1.53,
  2,       2,       2,       2,
  1.46,    1.46,    1.46,    1.46,
  1.37,    1.37,    1.37,    1.37,
  1.64,    1.64,    1.64,    1.64,
  1.95,    1.95,    1.95,    1.95,
  2.05,    2.05,    2.05,    2.05,
  1.79,    1.79,    1.79,    1.79,
  1.33,    1.33,    1.33,    1.33,
  1.65,    1.65,    1.65,    1.65,
  1.58,    1.58,    1.58,    1.58,
  1.97,    1.97,    1.97,    1.97,
  2,       2,       2,       2,
  2.05,    2.05,    2.05,    2.05,
  2.3,     2.3,     2.3,     2.3,
  2.24,    2.24,    2.24,    2.24,
  2.08,    2.08,    2.08,    2.08,
  1.79,    1.79,    1.79,    1.79,
  1.57,    1.57,    1.57,    1.57,
  1.95,    1.95,    1.95,    1.95,
  1.79,    1.79,    1.79,    1.79,
  1.76,    1.76,    1.76,    1.76,
  1.68,    1.68,    1.68,    1.68,
  1.6,     1.6,     1.6,     1.6,
  1.9,     1.9,     1.9,     1.9,
  1.76,    1.76,    1.76,    1.76,
  1.93,    1.93,    1.93,    1.93,
  1.89,    1.89,    1.89,    1.89,
  2.07,    2.07,    2.07,    2.07,
  2.43,    2.43,    2.43,    2.43,
  1.556,   1.556,   1.556,   1.556,
  2.85,    2.85,    2.85,    2.85,
  2.6,     2.6,     2.6,     2.6,
  2.61,    2.61,    2.61,    2.61,
  2.64,    2.64,    2.64,    2.64,
  3.04,    3.04,    3.04,    3.04,
  2.76,    2.76,    2.76,    2.76,
  2.83,    2.83,    2.83,    2.83,
  2.91,    2.91,    2.91,    2.91,
  3.02,    3.02,    3.02,    3.02,
  3.2,     3.2,     3.2,     3.2,
  2.97,    2.97,    2.97,    2.97,
  3.31,    3.31,    3.31,    3.31,
  3.62,    3.62,    3.62,    3.62,
  3.47,    3.47,    3.47,    3.47,
  3.75,    3.75,    3.75,    3.75,
  3.45,    3.45,    3.45,    3.45,
  3.79,    3.79,    3.79,    3.79,
  3.81,    3.81,    3.81,    3.81,
  3.83,    3.83,    3.83,    3.83,
  4.01,    4.01,    4.01,    4.01,
  3.98,    3.98,    3.98,    3.98,
  3.82,    3.82,    3.82,    3.82,
  3.85,    3.85,    3.85,    3.85,
  3.81,    3.81,    3.81,    3.81,
  3.7,     3.7,     3.7,     3.7,
  3.52,    3.52,    3.52,    3.52,
  3.67,    3.67,    3.67,    3.67,
  3.87,    3.87,    3.87,    3.87,
  3.7,     3.7,     3.7,     3.7,
  3.11,    3.11,    3.11,    3.11,
  3.08,    3.08,    3.08,    3.08,
  3.33,    3.33,    3.33,    3.33,
  3.41,    3.41,    3.41,    3.41,
  3.51,    3.51,    3.51,    3.51,
  3.21,    3.21,    3.21,    3.21,
  3.09,    3.09,    3.09,    3.09,
  3.28,    3.28,    3.28,    3.28,
  3.02,    3.02,    3.02,    3.02,
  3.2,     3.2,     3.2,     3.2,
  3.23,    3.23,    3.23,    3.23,
  3.24,    3.24,    3.24,    3.24,
  2.96,    2.96,    2.96,    2.96,
  2.87,    2.87,    2.87,    2.87,
  2.69,    2.69,    2.69,    2.69,
  2.09,    2.09,    2.09,    2.09,
  2.29,    2.29,    2.29,    2.29,
  2.56,    2.56,    2.56,    2.56,
  2.82,    2.82,    2.82,    2.82,
  3.19,    3.19,    3.19,    3.19,
  2.96,    2.96,    2.96,    2.96,
  2.94,    2.94,    2.94,    2.94,
  2.53,    2.53,    2.53,    2.53,
  2.29,    2.29,    2.29,    2.29,
  2.4,     2.4,     2.4,     2.4,
  2.74,    2.74,    2.74,    2.74,
  2.81,    2.81,    2.81,    2.81,
  2.52,    2.52,    2.52,    2.52,
  2.33,    2.33,    2.33,    2.33,
  2.65,    2.65,    2.65,    2.65,
  2.65,    2.65,    2.65,    2.65,
  2.45,    2.45,    2.45,    2.45,
  2.03,    2.03,    2.03,    2.03,
  2.24,    2.24,    2.24,    2.24,
  2.55,    2.55,    2.55,    2.55,
  2.43,    2.43,    2.43,    2.43,
  2.31,    2.31,    2.31,    2.31,
  2.65,    2.65,    2.65,    2.65,
  2.43,    2.43,    2.43,    2.43,
  2.46,    2.46,    2.46,    2.46,
  1.97,    1.97,    1.97,    1.97,
  2.13,    2.13,    2.13,    2.13,
  2.16,    2.16,    2.16,    2.16,
  1.93,    1.93,    1.93,    1.93,
  1.92,    1.92,    1.92,    1.92,
  2.51,    2.51,    2.51,    2.51,
  2.48,    2.48,    2.48,    2.48,
  2.65,    2.65,    2.65,    2.65,
  2.88,    2.88,    2.88,    2.88,
  2.63,    2.63,    2.63,    2.63,
  2.56,    2.56,    2.56,    2.56,
  2.52,    2.52,    2.52,    2.52,
  2.5,     2.5,     2.5,     2.5,
  2.56,    2.56,    2.56,    2.56,
  2.63,    2.63,    2.63,    2.63,
  2.36,    2.36,    2.36,    2.36,
  2.47,    2.47,    2.47,    2.47,
  2.01,    2.01,    2.01,    2.01,
  2.03,    2.03,    2.03,    2.03,
  2.24,    2.24,    2.24,    2.24,
  2.02,    2.02,    2.02,    2.02,
  2.29,    2.29,    2.29,    2.29,
  2.71,    2.71,    2.71,    2.71,
  2.13,    2.13,    2.13,    2.13,
  2.38,    2.38,    2.38,    2.38,
  2.21,    2.21,    2.21,    2.21,
  2.06,    2.06,    2.06,    2.06,
  1.77,    1.77,    1.77,    1.77,
  1.6,     1.6,     1.6,     1.6,
  0.96,    0.96,    0.96,    0.96,
  1.26,    1.26,    1.26,    1.26,
  1.92,    1.92,    1.92,    1.92,
  1.91,    1.91,    1.91,    1.91,
  1.37,    1.37,    1.37,    1.37,
  1.82,    1.82,    1.82,    1.82,
  1.84,    1.84,    1.84,    1.84,
  2.1,     2.1,     2.1,     2.1,
  1.84,    1.84,    1.84,    1.84,
  1.82,    1.82,    1.82,    1.82,
  1.8,     1.8,     1.8,     1.8,
  1.8,     1.8,     1.8,     1.8,
  1.5,     1.5,     1.5,     1.5,
  1.6,     1.6,     1.6,     1.6,
  1.22,    1.22,    1.22,    1.22,
  1.67,    1.67,    1.67,    1.67,
  1.62,    1.62,    1.62,    1.62,
  1.55,    1.55,    1.55,    1.55,
  1.64,    1.64,    1.64,    1.64,
  0.93,    0.93,    0.93,    0.93,
  0.98,    0.98,    0.98,    0.98,
  1.64,    1.64,    1.64,    1.64,
  1.53,    1.53,    1.53,    1.53,
  1.01,    1.01,    1.01,    1.01,
  1.77,    1.77,    1.77,    1.77,
  1.45,    1.45,    1.45,    1.45,
  2.05,    2.05,    2.05,    2.05,
  1.56,    1.56,    1.56,    1.56,
  1.61,    1.61,    1.61,    1.61,
  1.26,    1.26,    1.26,    1.26,
  1.09,    1.09,    1.09,    1.09,
  1.37,    1.37,    1.37,    1.37,
  1.09,    1.09,    1.09,    1.09,
  0.51,    0.51,    0.51,    0.51,
  0.41,    0.41,    0.41,    0.41,
  0.39,    0.39,    0.39,    0.39,
  0.68,    0.68,    0.68,    0.68,
  0.42,    0.42,    0.42,    0.42,
  0.43,    0.43,    0.43,    0.43,
  0.37,    0.37,    0.37,    0.37,
  0.25,    0.25,    0.25,    0.25,
  0.33,    0.33,    0.33,    0.33,
  0.46,    0.46,    0.46,    0.46,
  0.62,    0.62,    0.62,    0.62,
  0.99,    0.99,    0.99,    0.99,
  0.7,     0.7,     0.7,     0.7,
  0.46,    0.46,    0.46,    0.46,
  0.63,    0.63,    0.63,    0.63,
  0.86,    0.86,    0.86,    0.86,
  0.64,    0.64,    0.64,    0.64,
  0.74,    0.74,    0.74,    0.74,
  0.99,    0.99,    0.99,    0.99,
  1.12,    1.12,    1.12,    1.12,
  0.29,    0.29,    0.29,    0.29,
  0.59,    0.59,    0.59,    0.59,
  1.67,    1.67,    1.67,    1.67,
  1.35,    1.35,    1.35,    1.35,
  0.53,    0.53,    0.53,    0.53,
  0.69,    0.69,    0.69,    0.69,
  1.54,    1.54,    1.54,    1.54,
  1.36,    1.36,    1.36,    1.36,
  1.39,    1.39,    1.39,    1.39,
  1.27,    1.27,    1.27,    1.27,
  1.55,    1.55,    1.55,    1.55,
  1.76,    1.76,    1.76,    1.76,
  0.71,    0.71,    0.71,    0.71,
  0.42,    0.42,    0.42,    0.42,
  1.42,    1.42,    1.42,    1.42,
  0.9,     0.9,     0.9,     0.9,
  1.11,    1.11,    1.11,    1.11,
  1.46,    1.46,    1.46,    1.46,
  1.86,    1.86,    1.86,    1.86,
  1.28,    1.28,    1.28,    1.28,
  1.3,     1.3,     1.3,     1.3,
  1.51,    1.51,    1.51,    1.51,
  1.32,    1.32,    1.32,    1.32,
  1.55,    1.55,    1.55,    1.55,
  0.99,    0.99,    0.99,    0.99,
  1.61,    1.61,    1.61,    1.61,
  1.41,    1.41,    1.41,    1.41,
  1.58,    1.58,    1.58,    1.58,
  1.34,    1.34,    1.34,    1.34,
  1.39,    1.39,    1.39,    1.39,
  1.5,     1.5,     1.5,     1.5,
  0.86,    0.86,    0.86,    0.86,
  0.44,    0.44,    0.44,    0.44,
  0.65,    0.65,    0.65,    0.65,
  0.66,    0.66,    0.66,    0.66,
  0.81,    0.81,    0.81,    0.81,
  0.7,     0.7,     0.7,     0.7,
  0.94,    0.94,    0.94,    0.94,
  0.66,    0.66,    0.66,    0.66,
  0.29,    0.29,    0.29,    0.29,
  0.48,    0.48,    0.48,    0.48,
  1.09,    1.09,    1.09,    1.09,
  1.72,    1.72,    1.72,    1.72,
  1.79,    1.79,    1.79,    1.79,
  2.01,    2.01,    2.01,    2.01,
  2.37,    2.37,    2.37,    2.37,
  2.53,    2.53,    2.53,    2.53,
  1.54,    1.54,    1.54,    1.54,
  1.01,    1.01,    1.01,    1.01,
  1.38,    1.38,    1.38,    1.38,
  2.43,    2.43,    2.43,    2.43,
  2.1,     2.1,     2.1,     2.1,
  1.6,     1.6,     1.6,     1.6,
  1.33,    1.33,    1.33,    1.33,
  1.53,    1.53,    1.53,    1.53,
  1.15,    1.15,    1.15,    1.15,
  1.11,    1.11,    1.11,    1.11,
  1.58,    1.58,    1.58,    1.58,
  1.56,    1.56,    1.56,    1.56,
  1.85,    1.85,    1.85,    1.85,
  2.45,    2.45,    2.45,    2.45,
  2.1,     2.1,     2.1,     2.1,
  1.82,    1.82,    1.82,    1.82,
  0.79,    0.79,    0.79,    0.79,
  1.16,    1.16,    1.16,    1.16,
  1.26,    1.26,    1.26,    1.26,
  1.34,    1.34,    1.34,    1.34,
  1.51,    1.51,    1.51,    1.51,
  1.57,    1.57,    1.57,    1.57,
  1.54,    1.54,    1.54,    1.54,
  1.63,    1.63,    1.63,    1.63,
  1.68,    1.68,    1.68,    1.68,
  1.57,    1.57,    1.57,    1.57,
  1.36,    1.36,    1.36,    1.36,
  1.32,    1.32,    1.32,    1.32,
  1.91,    1.91,    1.91,    1.91,
  2.87,    2.87,    2.87,    2.87,
  2.51,    2.51,    2.51,    2.51,
  3.2,     3.2,     3.2,     3.2,
  2.83,    2.83,    2.83,    2.83,
  3.18,    3.18,    3.18,    3.18,
  3.41,    3.41,    3.41,    3.41,
  2.9,     2.9,     2.9,     2.9,
  2.76,    2.76,    2.76,    2.76,
  2.5,     2.5,     2.5,     2.5,
  1.3,     1.3,     1.3,     1.3,
  1.64,    1.64,    1.64,    1.64,
  1.68,    1.68,    1.68,    1.68,
  1.63,    1.63,    1.63,    1.63,
  1.69,    1.69,    1.69,    1.69,
  1.83,    1.83,    1.83,    1.83,
  2.02,    2.02,    2.02,    2.02,
  2.15,    2.15,    2.15,    2.15,
  2.24,    2.24,    2.24,    2.24,
  1.34,    1.34,    1.34,    1.34,
  0.43,    0.43,    0.43,    0.43,
  0.88,    0.88,    0.88,    0.88,
  1.57,    1.57,    1.57,    1.57,
  1.9,     1.9,     1.9,     1.9,
  1.39,    1.39,    1.39,    1.39,
  1.49,    1.49,    1.49,    1.49,
  1.48,    1.48,    1.48,    1.48,
  1.77,    1.77,    1.77,    1.77,
  1.73,    1.73,    1.73,    1.73,
  1.77,    1.77,    1.77,    1.77,
  1.8,     1.8,     1.8,     1.8,
  1.85,    1.85,    1.85,    1.85,
  1.79,    1.79,    1.79,    1.79,
  1.74,    1.74,    1.74,    1.74,
  1.66,    1.66,    1.66,    1.66,
  2.02,    2.02,    2.02,    2.02,
  1.88,    1.88,    1.88,    1.88,
  1.71,    1.71,    1.71,    1.71,
  1.75,    1.75,    1.75,    1.75,
  1.38,    1.38,    1.38,    1.38,
  1.24,    1.24,    1.24,    1.24,
  1.48,    1.48,    1.48,    1.48,
  1.57,    1.57,    1.57,    1.57,
  1.47,    1.47,    1.47,    1.47,
  1.66,    1.66,    1.66,    1.66,
  1.69,    1.69,    1.69,    1.69,
  1.24,    1.24,    1.24,    1.24,
  1.69,    1.69,    1.69,    1.69,
  2.1,     2.1,     2.1,     2.1,
  1,       1,       1,       1,
  1.69,    1.69,    1.69,    1.69,
  1.98,    1.98,    1.98,    1.98,
  1.43,    1.43,    1.43,    1.43,
  0.84,    0.84,    0.84,    0.84,
  1.18,    1.18,    1.18,    1.18,
  0.86,    0.86,    0.86,    0.86,
  1.07,    1.07,    1.07,    1.07,
  0.79,    0.79,    0.79,    0.79,
  0.68,    0.68,    0.68,    0.68,
  0.47,    0.47,    0.47,    0.47,
  1.11,    1.11,    1.11,    1.11,
  0.7,     0.7,     0.7,     0.7,
  0.81,    0.81,    0.81,    0.81,
  0.65,    0.65,    0.65,    0.65,
  1.41,    1.41,    1.41,    1.41,
  0.38,    0.38,    0.38,    0.38,
  0.54,    0.54,    0.54,    0.54,
  1.18,    1.18,    1.18,    1.18,
  0.82,    0.82,    0.82,    0.82,
  0.84,    0.84,    0.84,    0.84,
  1.53,    1.53,    1.53,    1.53,
  1.43,    1.43,    1.43,    1.43,
  1.49,    1.49,    1.49,    1.49,
  1.82,    1.82,    1.82,    1.82,
  1.71,    1.71,    1.71,    1.71,
  1.15,    1.15,    1.15,    1.15,
  0.74,    0.74,    0.74,    0.74,
  0.84,    0.84,    0.84,    0.84,
  1.27,    1.27,    1.27,    1.27,
  0.82,    0.82,    0.82,    0.82,
  1.35,    1.35,    1.35,    1.35,
  1.99,    1.99,    1.99,    1.99,
  0.63,    0.63,    0.63,    0.63,
  0.52,    0.52,    0.52,    0.52,
  0.47,    0.47,    0.47,    0.47,
  0.48,    0.48,    0.48,    0.48,
  0.43,    0.43,    0.43,    0.43,
  0.84,    0.84,    0.84,    0.84,
  0.73,    0.73,    0.73,    0.73,
  0.58,    0.58,    0.58,    0.58,
  0.57,    0.57,    0.57,    0.57,
  0.7,     0.7,     0.7,     0.7,
  0.91,    0.91,    0.91,    0.91,
  1.2,     1.2,     1.2,     1.2,
  1.13,    1.13,    1.13,    1.13,
  1.08,    1.08,    1.08,    1.08,
  1.57,    1.57,    1.57,    1.57,
  1.52,    1.52,    1.52,    1.52,
  1.1,     1.1,     1.1,     1.1,
  1.12,    1.12,    1.12,    1.12,
  1.18,    1.18,    1.18,    1.18,
  0.89,    0.89,    0.89,    0.89,
  1.11,    1.11,    1.11,    1.11,
  1.11,    1.11,    1.11,    1.11,
  1.15,    1.15,    1.15,    1.15,
  1.6,     1.6,     1.6,     1.6,
  1.79,    1.79,    1.79,    1.79,
  2.13,    2.13,    2.13,    2.13,
  1.74,    1.74,    1.74,    1.74,
  1.49,    1.49,    1.49,    1.49,
  1.55,    1.55,    1.55,    1.55,
  1.15,    1.15,    1.15,    1.15,
  1.5,     1.5,     1.5,     1.5,
  1.45,    1.45,    1.45,    1.45,
  1.16,    1.16,    1.16,    1.16,
  1.38,    1.38,    1.38,    1.38,
  1.6,     1.6,     1.6,     1.6,
  1.21,    1.21,    1.21,    1.21,
  0.98,    0.98,    0.98,    0.98,
  1.05,    1.05,    1.05,    1.05,
  1.29,    1.29,    1.29,    1.29,
  1.33,    1.33,    1.33,    1.33,
  1.8,     1.8,     1.8,     1.8,
  1.64,    1.64,    1.64,    1.64,
  1.65,    1.65,    1.65,    1.65,
  1.53,    1.53,    1.53,    1.53,
  1.15,    1.15,    1.15,    1.15,
  1.69,    1.69,    1.69,    1.69,
  1.58,    1.58,    1.58,    1.58,
  1.44,    1.44,    1.44,    1.44,
  1.25,    1.25,    1.25,    1.25,
  1.32,    1.32,    1.32,    1.32,
  0.97,    0.97,    0.97,    0.97,
  0.7,     0.7,     0.7,     0.7,
  0.75,    0.75,    0.75,    0.75,
  0.96,    0.96,    0.96,    0.96,
  1.49,    1.49,    1.49,    1.49,
  1.32,    1.32,    1.32,    1.32,
  1.75,    1.75,    1.75,    1.75,
  1.3,     1.3,     1.3,     1.3,
  2.15,    2.15,    2.15,    2.15,
  1.97,    1.97,    1.97,    1.97,
  1.88,    1.88,    1.88,    1.88,
  1.85,    1.85,    1.85,    1.85,
  1.63,    1.63,    1.63,    1.63,
  2.09,    2.09,    2.09,    2.09,
  2.06,    2.06,    2.06,    2.06,
  1.6,     1.6,     1.6,     1.6,
  1.24,    1.24,    1.24,    1.24,
  1.49,    1.49,    1.49,    1.49,
  1,       1,       1,       1,
  0.87,    0.87,    0.87,    0.87,
  0.61,    0.61,    0.61,    0.61,
  0.78,    0.78,    0.78,    0.78,
  0.64,    0.64,    0.64,    0.64,
  0.31,    0.31,    0.31,    0.31,
  0.11,    0.11,    0.11,    0.11,
  1.19,    1.19,    1.19,    1.19,
  1.08,    1.08,    1.08,    1.08,
  0.9,     0.9,     0.9,     0.9,
  0.93,    0.93,    0.93,    0.93,
  1.24,    1.24,    1.24,    1.24,
  1.2,     1.2,     1.2,     1.2,
  0.71,    0.71,    0.71,    0.71,
  0.63,    0.63,    0.63,    0.63,
  0.9,     0.9,     0.9,     0.9,
  0.84,    0.84,    0.84,    0.84,
  0.64,    0.64,    0.64,    0.64,
  0.44,    0.44,    0.44,    0.44,
  0.72,    0.72,    0.72,    0.72,
  0.56,    0.56,    0.56,    0.56,
  0.28,    0.28,    0.28,    0.28,
  0.26,    0.26,    0.26,    0.26,
  0.21,    0.21,    0.21,    0.21,
  0.17,    0.17,    0.17,    0.17,
  0.03,    0.03,    0.03,    0.03,
  0.35,    0.35,    0.35,    0.35,
  0.42,    0.42,    0.42,    0.42,
  0.72,    0.72,    0.72,    0.72,
  0.46,    0.46,    0.46,    0.46,
  0.69,    0.69,    0.69,    0.69,
  0.57,    0.57,    0.57,    0.57,
  0.77,    0.77,    0.77,    0.77,
  0.87,    0.87,    0.87,    0.87,
  0.38,    0.38,    0.38,    0.38,
  0.36,    0.36,    0.36,    0.36,
  0.98,    0.98,    0.98,    0.98,
  0.66,    0.66,    0.66,    0.66,
  0.91,    0.91,    0.91,    0.91,
  1.29,    1.29,    1.29,    1.29,
  1.24,    1.24,    1.24,    1.24,
  1.02,    1.02,    1.02,    1.02,
  0.89,    0.89,    0.89,    0.89,
  1.14,    1.14,    1.14,    1.14,
  1.14,    1.14,    1.14,    1.14,
  1.09,    1.09,    1.09,    1.09,
  0.47,    0.47,    0.47,    0.47,
  0.49,    0.49,    0.49,    0.49,
  0.26,    0.26,    0.26,    0.26,
  0.54,    0.54,    0.54,    0.54,
  0.99,    0.99,    0.99,    0.99,
  1.03,    1.03,    1.03,    1.03,
  0.87,    0.87,    0.87,    0.87,
  0.88,    0.88,    0.88,    0.88,
  0.72,    0.72,    0.72,    0.72,
  0.84,    0.84,    0.84,    0.84,
  1.05,    1.05,    1.05,    1.05,
  1.13,    1.13,    1.13,    1.13,
  1.15,    1.15,    1.15,    1.15,
  1.05,    1.05,    1.05,    1.05,
  1.12,    1.12,    1.12,    1.12,
  0.66,    0.66,    0.66,    0.66,
  0.69,    0.69,    0.69,    0.69,
  0.94,    0.94,    0.94,    0.94,
  1.08,    1.08,    1.08,    1.08,
  1.22,    1.22,    1.22,    1.22,
  1,       1,       1,       1,
  1.13,    1.13,    1.13,    1.13,
  1.19,    1.19,    1.19,    1.19,
  1.38,    1.38,    1.38,    1.38,
  1.51,    1.51,    1.51,    1.51,
  1.15,    1.15,    1.15,    1.15,
  1.27,    1.27,    1.27,    1.27,
  1.08,    1.08,    1.08,    1.08,
  1.17,    1.17,    1.17,    1.17,
  1.24,    1.24,    1.24,    1.24,
  1.37,    1.37,    1.37,    1.37,
  1.1,     1.1,     1.1,     1.1,
  1.06,    1.06,    1.06,    1.06,
  1.58,    1.58,    1.58,    1.58,
  1.44,    1.44,    1.44,    1.44,
  1.73,    1.73,    1.73,    1.73,
  1.99,    1.99,    1.99,    1.99,
  1.95,    1.95,    1.95,    1.95,
  2.18,    2.18,    2.18,    2.18,
  2.27,    2.27,    2.27,    2.27,
  2.3,     2.3,     2.3,     2.3,
  2.34,    2.34,    2.34,    2.34,
  2.01,    2.01,    2.01,    2.01,
  1.6,     1.6,     1.6,     1.6,
  1.69,    1.69,    1.69,    1.69,
  1.25,    1.25,    1.25,    1.25,
  1.19,    1.19,    1.19,    1.19,
  1.64,    1.64,    1.64,    1.64,
  1.86,    1.86,    1.86,    1.86,
  1.5,     1.5,     1.5,     1.5,
  1.78,    1.78,    1.78,    1.78,
  1.85,    1.85,    1.85,    1.85,
  1.75,    1.75,    1.75,    1.75,
  1.62,    1.62,    1.62,    1.62,
  1.33,    1.33,    1.33,    1.33,
  1.96,    1.96,    1.96,    1.96,
  2.21,    2.21,    2.21,    2.21,
  1.8,     1.8,     1.8,     1.8,
  2.18,    2.18,    2.18,    2.18,
  1.44,    1.44,    1.44,    1.44,
  1.21,    1.21,    1.21,    1.21,
  1.28,    1.28,    1.28,    1.28,
  1.66,    1.66,    1.66,    1.66,
  1.41,    1.41,    1.41,    1.41,
  1.67,    1.67,    1.67,    1.67,
  1.56,    1.56,    1.56,    1.56,
  1.89,    1.89,    1.89,    1.89,
  1.74,    1.74,    1.74,    1.74,
  1.7,     1.7,     1.7,     1.7,
  1.52,    1.52,    1.52,    1.52,
  1.29,    1.29,    1.29,    1.29,
  1.3,     1.3,     1.3,     1.3,
  1.47,    1.47,    1.47,    1.47,
  1.38,    1.38,    1.38,    1.38,
  1.08,    1.08,    1.08,    1.08,
  0.57,    0.57,    0.57,    0.57,
  0.99,    0.99,    0.99,    0.99,
  0.8,     0.8,     0.8,     0.8,
  1.34,    1.34,    1.34,    1.34,
  1.01,    1.01,    1.01,    1.01,
  0.66,    0.66,    0.66,    0.66,
  1.03,    1.03,    1.03,    1.03,
  1.57,    1.57,    1.57,    1.57,
  1.21,    1.21,    1.21,    1.21,
  0.98,    0.98,    0.98,    0.98,
  1.56,    1.56,    1.56,    1.56,
  1.5,     1.5,     1.5,     1.5,
  1.19,    1.19,    1.19,    1.19,
  0.87,    0.87,    0.87,    0.87,
  0.71,    0.71,    0.71,    0.71,
  0.99,    0.99,    0.99,    0.99,
  1.41,    1.41,    1.41,    1.41,
  1.36,    1.36,    1.36,    1.36,
  1.43,    1.43,    1.43,    1.43,
  1.49,    1.49,    1.49,    1.49,
  1.31,    1.31,    1.31,    1.31,
  1.52,    1.52,    1.52,    1.52,
  1.52,    1.52,    1.52,    1.52,
  0.86,    0.86,    0.86,    0.86,
  1.33,    1.33,    1.33,    1.33,
  2.04,    2.04,    2.04,    2.04,
  2.25,    2.25,    2.25,    2.25,
  1.88,    1.88,    1.88,    1.88,
  2.32,    2.32,    2.32,    2.32,
  2.14,    2.14,    2.14,    2.14,
  2.49,    2.49,    2.49,    2.49,
  1.73,    1.73,    1.73,    1.73,
  2.29,    2.29,    2.29,    2.29,
  2.13,    2.13,    2.13,    2.13,
  2.07,    2.07,    2.07,    2.07,
  1.66,    1.66,    1.66,    1.66,
  1.8,     1.8,     1.8,     1.8,
  1.3,     1.3,     1.3,     1.3,
  1.31,    1.31,    1.31,    1.31,
  1.55,    1.55,    1.55,    1.55,
  1.47,    1.47,    1.47,    1.47,
  1.79,    1.79,    1.79,    1.79,
  1.72,    1.72,    1.72,    1.72,
  1.95,    1.95,    1.95,    1.95,
  2.09,    2.09,    2.09,    2.09,
  2.21,    2.21,    2.21,    2.21,
  2.16,    2.16,    2.16,    2.16,
  2.46,    2.46,    2.46,    2.46,
  2.24,    2.24,    2.24,    2.24,
  2.14,    2.14,    2.14,    2.14,
  1.97,    1.97,    1.97,    1.97,
  2.23,    2.23,    2.23,    2.23,
  2.32,    2.32,    2.32,    2.32,
  2.3,     2.3,     2.3,     2.3,
  2.36,    2.36,    2.36,    2.36,
  2.54,    2.54,    2.54,    2.54,
  2.51,    2.51,    2.51,    2.51,
  2.29,    2.29,    2.29,    2.29,
  2.24,    2.24,    2.24,    2.24,
  2.33,    2.33,    2.33,    2.33,
  2.07,    2.07,    2.07,    2.07,
  2.24,    2.24,    2.24,    2.24,
  2.12,    2.12,    2.12,    2.12,
  2.06,    2.06,    2.06,    2.06,
  1.95,    1.95,    1.95,    1.95,
  2.17,    2.17,    2.17,    2.17,
  2.52,    2.52,    2.52,    2.52,
  2.57,    2.57,    2.57,    2.57,
  2.23,    2.23,    2.23,    2.23,
  1.92,    1.92,    1.92,    1.92,
  2.07,    2.07,    2.07,    2.07,
  2.33,    2.33,    2.33,    2.33,
  2.31,    2.31,    2.31,    2.31,
  1.89,    1.89,    1.89,    1.89,
  2.04,    2.04,    2.04,    2.04,
  2.7,     2.7,     2.7,     2.7,
  2.32,    2.32,    2.32,    2.32,
  2.78,    2.78,    2.78,    2.78,
  2.79,    2.79,    2.79,    2.79,
  2.09,    2.09,    2.09,    2.09,
  2.87,    2.87,    2.87,    2.87,
  2.76,    2.76,    2.76,    2.76,
  2.28,    2.28,    2.28,    2.28,
  2.2,     2.2,     2.2,     2.2,
  2.11,    2.11,    2.11,    2.11,
  2.27,    2.27,    2.27,    2.27,
  2.07,    2.07,    2.07,    2.07,
  2.18,    2.18,    2.18,    2.18,
  2.06,    2.06,    2.06,    2.06,
  1.98,    1.98,    1.98,    1.98,
  1.72,    1.72,    1.72,    1.72,
  1.88,    1.88,    1.88,    1.88,
  1.98,    1.98,    1.98,    1.98,
  1.92,    1.92,    1.92,    1.92,
  1.63,    1.63,    1.63,    1.63,
  1.63,    1.63,    1.63,    1.63,
  1.54,    1.54,    1.54,    1.54,
  1.41,    1.41,    1.41,    1.41,
  1.48,    1.48,    1.48,    1.48,
  1.47,    1.47,    1.47,    1.47,
  1.45,    1.45,    1.45,    1.45,
  1.14,    1.14,    1.14,    1.14,
  1.22,    1.22,    1.22,    1.22,
  1.25,    1.25,    1.25,    1.25,
  1.24,    1.24,    1.24,    1.24,
  0.97,    0.97,    0.97,    0.97,
  0.93,    0.93,    0.93,    0.93,
  0.93,    0.93,    0.93,    0.93,
  1.46,    1.46,    1.46,    1.46,
  1.16,    1.16,    1.16,    1.16,
  1.63,    1.63,    1.63,    1.63,
  1.64,    1.64,    1.64,    1.64,
  1.81,    1.81,    1.81,    1.81,
  1.05,    1.05,    1.05,    1.05,
  0.82,    0.82,    0.82,    0.82,
  1.11,    1.11,    1.11,    1.11,
  0.46,    0.46,    0.46,    0.46,
  0.76,    0.76,    0.76,    0.76,
  0.94,    0.94,    0.94,    0.94,
  0.88,    0.88,    0.88,    0.88,
  1.01,    1.01,    1.01,    1.01,
  1.11,    1.11,    1.11,    1.11,
  1.68,    1.68,    1.68,    1.68,
  1.45,    1.45,    1.45,    1.45,
  1.45,    1.45,    1.45,    1.45,
  1.57,    1.57,    1.57,    1.57,
  1.91,    1.91,    1.91,    1.91,
  1.99,    1.99,    1.99,    1.99,
  1.65,    1.65,    1.65,    1.65,
  1.87,    1.87,    1.87,    1.87,
  2.54,    2.54,    2.54,    2.54,
  1.93,    1.93,    1.93,    1.93,
  2.79,    2.79,    2.79,    2.79,
  2.92,    2.92,    2.92,    2.92,
  2.77,    2.77,    2.77,    2.77,
  2.72,    2.72,    2.72,    2.72,
  2.87,    2.87,    2.87,    2.87,
  2.68,    2.68,    2.68,    2.68,
  2.44,    2.44,    2.44,    2.44,
  3.21,    3.21,    3.21,    3.21,
  3.18,    3.18,    3.18,    3.18,
  3.17,    3.17,    3.17,    3.17,
  3.38,    3.38,    3.38,    3.38,
  3.45,    3.45,    3.45,    3.45,
  3.34,    3.34,    3.34,    3.34,
  3.25,    3.25,    3.25,    3.25,
  3.36,    3.36,    3.36,    3.36,
  3.26,    3.26,    3.26,    3.26,
  3.62,    3.62,    3.62,    3.62,
  3.94,    3.94,    3.94,    3.94,
  4.21,    4.21,    4.21,    4.21,
  4.33,    4.33,    4.33,    4.33,
  4.54,    4.54,    4.54,    4.54,
  4.46,    4.46,    4.46,    4.46,
  4.34,    4.34,    4.34,    4.34,
  3.91,    3.91,    3.91,    3.91,
  4.14,    4.14,    4.14,    4.14,
  4.18,    4.18,    4.18,    4.18,
  4.36,    4.36,    4.36,    4.36,
  4.94,    4.94,    4.94,    4.94,
  4.73,    4.73,    4.73,    4.73,
  4.76,    4.76,    4.76,    4.76,
  4.59,    4.59,    4.59,    4.59,
  4.11,    4.11,    4.11,    4.11,
  4.29,    4.29,    4.29,    4.29,
  4.85,    4.85,    4.85,    4.85,
  4.59,    4.59,    4.59,    4.59,
  4.71,    4.71,    4.71,    4.71,
  4.52,    4.52,    4.52,    4.52,
  5.34,    5.34,    5.34,    5.34,
  5.28,    5.28,    5.28,    5.28,
  5.2,     5.2,     5.2,     5.2,
  4.9,     4.9,     4.9,     4.9,
  5.26,    5.26,    5.26,    5.26,
  4.94,    4.94,    4.94,    4.94,
  5.5,     5.5,     5.5,     5.5,
  5.21,    5.21,    5.21,    5.21,
  5.44,    5.44,    5.44,    5.44,
  5.66,    5.66,    5.66,    5.66,
  5.57,    5.57,    5.57,    5.57,
  5.62,    5.62,    5.62,    5.62,
  5.41,    5.41,    5.41,    5.41,
  5.78,    5.78,    5.78,    5.78,
  5.79,    5.79,    5.79,    5.79,
  5.25,    5.25,    5.25,    5.25,
  5.3,     5.3,     5.3,     5.3,
  5.28,    5.28,    5.28,    5.28,
  5.46,    5.46,    5.46,    5.46,
  5.35,    5.35,    5.35,    5.35,
  4.85,    4.85,    4.85,    4.85,
  4.26,    4.26,    4.26,    4.26,
  4.37,    4.37,    4.37,    4.37,
  4.56,    4.56,    4.56,    4.56,
  2.99,    2.99,    2.99,    2.99,
  2.57,    2.57,    2.57,    2.57,
  2.54,    2.54,    2.54,    2.54,
  2.37,    2.37,    2.37,    2.37,
  3.17,    3.17,    3.17,    3.17,
  2.23,    2.23,    2.23,    2.23,
  1.83,    1.83,    1.83,    1.83,
  1.16,    1.16,    1.16,    1.16,
  1.32,    1.32,    1.32,    1.32,
  1.88,    1.88,    1.88,    1.88,
  2.38,    2.38,    2.38,    2.38,
  2.12,    2.12,    2.12,    2.12,
  1.89,    1.89,    1.89,    1.89,
  2.02,    2.02,    2.02,    2.02,
  1.46,    1.46,    1.46,    1.46,
  1.87,    1.87,    1.87,    1.87,
  2.14,    2.14,    2.14,    2.14,
  1.94,    1.94,    1.94,    1.94,
  1.7,     1.7,     1.7,     1.7,
  1.74,    1.74,    1.74,    1.74,
  1.64,    1.64,    1.64,    1.64,
  1.78,    1.78,    1.78,    1.78,
  1.78,    1.78,    1.78,    1.78,
  2.35,    2.35,    2.35,    2.35,
  1.99,    1.99,    1.99,    1.99,
  1.78,    1.78,    1.78,    1.78,
  1.71,    1.71,    1.71,    1.71,
  2.27,    2.27,    2.27,    2.27,
  3.07,    3.07,    3.07,    3.07,
  3.09,    3.09,    3.09,    3.09,
  2.93,    2.93,    2.93,    2.93,
  2.64,    2.64,    2.64,    2.64,
  2.72,    2.72,    2.72,    2.72,
  2.31,    2.31,    2.31,    2.31,
  1.77,    1.77,    1.77,    1.77,
  1.44,    1.44,    1.44,    1.44,
  1.44,    1.44,    1.44,    1.44,
  2.08,    2.08,    2.08,    2.08,
  2.18,    2.18,    2.18,    2.18,
  2.27,    2.27,    2.27,    2.27,
  2.49,    2.49,    2.49,    2.49,
  2.49,    2.49,    2.49,    2.49,
  2.48,    2.48,    2.48,    2.48,
  2.28,    2.28,    2.28,    2.28,
  2.15,    2.15,    2.15,    2.15,
  2.24,    2.24,    2.24,    2.24,
  2.32,    2.32,    2.32,    2.32,
  2.34,    2.34,    2.34,    2.34,
  2.26,    2.26,    2.26,    2.26,
  2.41,    2.41,    2.41,    2.41,
  2.42,    2.42,    2.42,    2.42,
  2.46,    2.46,    2.46,    2.46,
  2.27,    2.27,    2.27,    2.27,
  2.26,    2.26,    2.26,    2.26,
  2.24,    2.24,    2.24,    2.24,
  2.25,    2.25,    2.25,    2.25,
  2.39,    2.39,    2.39,    2.39,
  2.54,    2.54,    2.54,    2.54,
  2.56,    2.56,    2.56,    2.56,
  2.29,    2.29,    2.29,    2.29,
  2.42,    2.42,    2.42,    2.42,
  2.07,    2.07,    2.07,    2.07,
  2.95,    2.95,    2.95,    2.95,
  3.01,    3.01,    3.01,    3.01,
  3.07,    3.07,    3.07,    3.07,
  3.17,    3.17,    3.17,    3.17,
  3.31,    3.31,    3.31,    3.31,
  3.64,    3.64,    3.64,    3.64,
  3.97,    3.97,    3.97,    3.97,
  3.33,    3.33,    3.33,    3.33,
  3.66,    3.66,    3.66,    3.66,
  3.59,    3.59,    3.59,    3.59,
  3.59,    3.59,    3.59,    3.59,
  3.73,    3.73,    3.73,    3.73,
  3.75,    3.75,    3.75,    3.75,
  3.67,    3.67,    3.67,    3.67,
  3.72,    3.72,    3.72,    3.72,
  3.76,    3.76,    3.76,    3.76,
  4.28,    4.28,    4.28,    4.28,
  3.9,     3.9,     3.9,     3.9,
  3.59,    3.59,    3.59,    3.59,
  3.68,    3.68,    3.68,    3.68,
  3.48,    3.48,    3.48,    3.48,
  3.53,    3.53,    3.53,    3.53,
  3.38,    3.38,    3.38,    3.38,
  3.38,    3.38,    3.38,    3.38,
  3.99,    3.99,    3.99,    3.99,
  3.84,    3.84,    3.84,    3.84,
  4.15,    4.15,    4.15,    4.15,
  3.94,    3.94,    3.94,    3.94,
  3.87,    3.87,    3.87,    3.87,
  3.96,    3.96,    3.96,    3.96,
  3.8,     3.8,     3.8,     3.8,
  4.22,    4.22,    4.22,    4.22,
  3.75,    3.75,    3.75,    3.75,
  3.94,    3.94,    3.94,    3.94,
  3.65,    3.65,    3.65,    3.65,
  4.3,     4.3,     4.3,     4.3,
  4.32,    4.32,    4.32,    4.32,
  4.02,    4.02,    4.02,    4.02,
  3.95,    3.95,    3.95,    3.95,
  3.97,    3.97,    3.97,    3.97,
  3.77,    3.77,    3.77,    3.77,
  4,       4,       4,       4,
  3.82,    3.82,    3.82,    3.82,
  3.77,    3.77,    3.77,    3.77,
  4.08,    4.08,    4.08,    4.08,
  3.66,    3.66,    3.66,    3.66,
  3.94,    3.94,    3.94,    3.94,
  3.72,    3.72,    3.72,    3.72,
  3.78,    3.78,    3.78,    3.78,
  3.27,    3.27,    3.27,    3.27,
  3.44,    3.44,    3.44,    3.44,
  3.91,    3.91,    3.91,    3.91,
  3.76,    3.76,    3.76,    3.76,
  3.79,    3.79,    3.79,    3.79,
  3.85,    3.85,    3.85,    3.85,
  3.72,    3.72,    3.72,    3.72,
  3.84,    3.84,    3.84,    3.84,
  3.79,    3.79,    3.79,    3.79,
  4.09,    4.09,    4.09,    4.09,
  3.76,    3.76,    3.76,    3.76,
  3.12,    3.12,    3.12,    3.12,
  3.79,    3.79,    3.79,    3.79,
  3.8,     3.8,     3.8,     3.8,
  3.82,    3.82,    3.82,    3.82,
  3.42,    3.42,    3.42,    3.42,
  3.7,     3.7,     3.7,     3.7,
  3.15,    3.15,    3.15,    3.15,
  3.17,    3.17,    3.17,    3.17,
  3.35,    3.35,    3.35,    3.35,
  3.36,    3.36,    3.36,    3.36,
  3.02,    3.02,    3.02,    3.02,
  2.99,    2.99,    2.99,    2.99,
  3.09,    3.09,    3.09,    3.09,
  2.7,     2.7,     2.7,     2.7,
  3.08,    3.08,    3.08,    3.08,
  2.15,    2.15,    2.15,    2.15,
  1.13,    1.13,    1.13,    1.13,
  1.39,    1.39,    1.39,    1.39,
  1.51,    1.51,    1.51,    1.51,
  1.89,    1.89,    1.89,    1.89,
  1.43,    1.43,    1.43,    1.43,
  1.6,     1.6,     1.6,     1.6,
  1.38,    1.38,    1.38,    1.38,
  1.77,    1.77,    1.77,    1.77,
  1.55,    1.55,    1.55,    1.55,
  1,       1,       1,       1,
  1.66,    1.66,    1.66,    1.66,
  1.61,    1.61,    1.61,    1.61,
  1.1,     1.1,     1.1,     1.1,
  1.11,    1.11,    1.11,    1.11,
  1.12,    1.12,    1.12,    1.12,
  1.18,    1.18,    1.18,    1.18,
  0.46,    0.46,    0.46,    0.46,
  0.63,    0.63,    0.63,    0.63,
  0.83,    0.83,    0.83,    0.83,
  1.21,    1.21,    1.21,    1.21,
  1.11,    1.11,    1.11,    1.11,
  1.05,    1.05,    1.05,    1.05,
  1.18,    1.18,    1.18,    1.18,
  1.2,     1.2,     1.2,     1.2,
  0.91,    0.91,    0.91,    0.91,
  1.62,    1.62,    1.62,    1.62,
  1.86,    1.86,    1.86,    1.86,
  1.03,    1.03,    1.03,    1.03,
  1.17,    1.17,    1.17,    1.17,
  1.67,    1.67,    1.67,    1.67,
  1.18,    1.18,    1.18,    1.18,
  1.7,     1.7,     1.7,     1.7,
  1.55,    1.55,    1.55,    1.55,
  1.95,    1.95,    1.95,    1.95,
  1.49,    1.49,    1.49,    1.49,
  1.58,    1.58,    1.58,    1.58,
  2.05,    2.05,    2.05,    2.05,
  1.88,    1.88,    1.88,    1.88,
  1.55,    1.55,    1.55,    1.55,
  1.92,    1.92,    1.92,    1.92,
  1.85,    1.85,    1.85,    1.85,
  1.84,    1.84,    1.84,    1.84,
  1.85,    1.85,    1.85,    1.85,
  1.91,    1.91,    1.91,    1.91,
  1.79,    1.79,    1.79,    1.79,
  2.15,    2.15,    2.15,    2.15,
  1.88,    1.88,    1.88,    1.88,
  1.91,    1.91,    1.91,    1.91,
  1.81,    1.81,    1.81,    1.81,
  1.89,    1.89,    1.89,    1.89,
  2.1,     2.1,     2.1,     2.1,
  1.78,    1.78,    1.78,    1.78,
  2.01,    2.01,    2.01,    2.01,
  2.33,    2.33,    2.33,    2.33,
  1.96,    1.96,    1.96,    1.96,
  2.02,    2.02,    2.02,    2.02,
  1.95,    1.95,    1.95,    1.95,
  1.68,    1.68,    1.68,    1.68,
  2.04,    2.04,    2.04,    2.04,
  2.4,     2.4,     2.4,     2.4,
  2.79,    2.79,    2.79,    2.79,
  2.84,    2.84,    2.84,    2.84,
  2.76,    2.76,    2.76,    2.76,
  2.97,    2.97,    2.97,    2.97,
  3.83,    3.83,    3.83,    3.83,
  4.13,    4.13,    4.13,    4.13,
  3.46,    3.46,    3.46,    3.46,
  3.48,    3.48,    3.48,    3.48,
  4.04,    4.04,    4.04,    4.04,
  3.84,    3.84,    3.84,    3.84,
  3.28,    3.28,    3.28,    3.28,
  2.73,    2.73,    2.73,    2.73,
  2.91,    2.91,    2.91,    2.91,
  3.16,    3.16,    3.16,    3.16,
  3.05,    3.05,    3.05,    3.05,
  3.5,     3.5,     3.5,     3.5,
  3.8,     3.8,     3.8,     3.8,
  3.86,    3.86,    3.86,    3.86,
  4.05,    4.05,    4.05,    4.05,
  3.73,    3.73,    3.73,    3.73,
  3.57,    3.57,    3.57,    3.57,
  3.72,    3.72,    3.72,    3.72,
  4.62,    4.62,    4.62,    4.62,
  4.87,    4.87,    4.87,    4.87,
  4.39,    4.39,    4.39,    4.39,
  5.1,     5.1,     5.1,     5.1,
  4.03,    4.03,    4.03,    4.03,
  3.1,     3.1,     3.1,     3.1,
  3.02,    3.02,    3.02,    3.02,
  3.22,    3.22,    3.22,    3.22,
  2.56,    2.56,    2.56,    2.56,
  2.23,    2.23,    2.23,    2.23,
  2.37,    2.37,    2.37,    2.37,
  2.05,    2.05,    2.05,    2.05,
  2.06,    2.06,    2.06,    2.06,
  2.12,    2.12,    2.12,    2.12,
  2.45,    2.45,    2.45,    2.45,
  2.59,    2.59,    2.59,    2.59,
  2.8,     2.8,     2.8,     2.8,
  3.19,    3.19,    3.19,    3.19,
  3.23,    3.23,    3.23,    3.23,
  2.88,    2.88,    2.88,    2.88,
  3.14,    3.14,    3.14,    3.14,
  3.4,     3.4,     3.4,     3.4,
  3.04,    3.04,    3.04,    3.04,
  2.86,    2.86,    2.86,    2.86,
  2.79,    2.79,    2.79,    2.79,
  2.73,    2.73,    2.73,    2.73,
  3.07,    3.07,    3.07,    3.07,
  3.15,    3.15,    3.15,    3.15,
  3.64,    3.64,    3.64,    3.64,
  3.12,    3.12,    3.12,    3.12,
  3.17,    3.17,    3.17,    3.17,
  2.92,    2.92,    2.92,    2.92,
  3.14,    3.14,    3.14,    3.14,
  3.59,    3.59,    3.59,    3.59,
  3.44,    3.44,    3.44,    3.44,
  3.42,    3.42,    3.42,    3.42,
  3.78,    3.78,    3.78,    3.78,
  3.81,    3.81,    3.81,    3.81,
  4.63,    4.63,    4.63,    4.63,
  4.15,    4.15,    4.15,    4.15,
  4.34,    4.34,    4.34,    4.34,
  4.6,     4.6,     4.6,     4.6,
  4.95,    4.95,    4.95,    4.95,
  5.1,     5.1,     5.1,     5.1,
  5.49,    5.49,    5.49,    5.49,
  5.44,    5.44,    5.44,    5.44,
  4.96,    4.96,    4.96,    4.96,
  5.55,    5.55,    5.55,    5.55,
  5.47,    5.47,    5.47,    5.47,
  5.63,    5.63,    5.63,    5.63,
  5.66,    5.66,    5.66,    5.66,
  5.18,    5.18,    5.18,    5.18,
  5.2,     5.2,     5.2,     5.2,
  5.08,    5.08,    5.08,    5.08,
  5.42,    5.42,    5.42,    5.42,
  5.4,     5.4,     5.4,     5.4,
  5.85,    5.85,    5.85,    5.85,
  5.23,    5.23,    5.23,    5.23,
  5.91,    5.91,    5.91,    5.91,
  5.99,    5.99,    5.99,    5.99,
  5.26,    5.26,    5.26,    5.26,
  5.43,    5.43,    5.43,    5.43,
  5.12,    5.12,    5.12,    5.12,
  4.95,    4.95,    4.95,    4.95,
  4.55,    4.55,    4.55,    4.55,
  4.72,    4.72,    4.72,    4.72,
  5.51,    5.51,    5.51,    5.51,
  5.48,    5.48,    5.48,    5.48,
  5.63,    5.63,    5.63,    5.63,
  5.63,    5.63,    5.63,    5.63,
  5.59,    5.59,    5.59,    5.59,
  5.51,    5.51,    5.51,    5.51,
  5.2,     5.2,     5.2,     5.2,
  5.56,    5.56,    5.56,    5.56,
  4.9,     4.9,     4.9,     4.9,
  4.3,     4.3,     4.3,     4.3,
  4.2,     4.2,     4.2,     4.2,
  3.84,    3.84,    3.84,    3.84,
  4.01,    4.01,    4.01,    4.01,
  4.34,    4.34,    4.34,    4.34,
  4.18,    4.18,    4.18,    4.18,
  3.62,    3.62,    3.62,    3.62,
  3.91,    3.91,    3.91,    3.91,
  3.83,    3.83,    3.83,    3.83,
  3.8,     3.8,     3.8,     3.8,
  3.48,    3.48,    3.48,    3.48,
  3.89,    3.89,    3.89,    3.89,
  4.41,    4.41,    4.41,    4.41,
  5.04,    5.04,    5.04,    5.04,
  4.99,    4.99,    4.99,    4.99,
  4.92,    4.92,    4.92,    4.92,
  4.86,    4.86,    4.86,    4.86,
  5.41,    5.41,    5.41,    5.41,
  5.71,    5.71,    5.71,    5.71,
  5.57,    5.57,    5.57,    5.57,
  5.45,    5.45,    5.45,    5.45,
  5.34,    5.34,    5.34,    5.34,
  5.73,    5.73,    5.73,    5.73,
  5.46,    5.46,    5.46,    5.46,
  5.38,    5.38,    5.38,    5.38,
  5.53,    5.53,    5.53,    5.53,
  5.11,    5.11,    5.11,    5.11,
  4.87,    4.87,    4.87,    4.87,
  4.57,    4.57,    4.57,    4.57,
  4.34,    4.34,    4.34,    4.34,
  4.08,    4.08,    4.08,    4.08,
  3.85,    3.85,    3.85,    3.85,
  3.16,    3.16,    3.16,    3.16,
  3.46,    3.46,    3.46,    3.46,
  3.39,    3.39,    3.39,    3.39,
  4.24,    4.24,    4.24,    4.24,
  4.45,    4.45,    4.45,    4.45,
  3.81,    3.81,    3.81,    3.81,
  3.42,    3.42,    3.42,    3.42,
  3.5,     3.5,     3.5,     3.5,
  3.02,    3.02,    3.02,    3.02,
  2.95,    2.95,    2.95,    2.95,
  3.28,    3.28,    3.28,    3.28,
  3.27,    3.27,    3.27,    3.27,
  4.11,    4.11,    4.11,    4.11,
  3.82,    3.82,    3.82,    3.82,
  3.2,     3.2,     3.2,     3.2,
  3.26,    3.26,    3.26,    3.26,
  3.57,    3.57,    3.57,    3.57,
  3.55,    3.55,    3.55,    3.55,
  4.03,    4.03,    4.03,    4.03,
  4.49,    4.49,    4.49,    4.49,
  5.11,    5.11,    5.11,    5.11,
  4.26,    4.26,    4.26,    4.26,
  3.99,    3.99,    3.99,    3.99,
  4.12,    4.12,    4.12,    4.12,
  4.37,    4.37,    4.37,    4.37,
  4.36,    4.36,    4.36,    4.36,
  4.7,     4.7,     4.7,     4.7,
  4.53,    4.53,    4.53,    4.53,
  4.39,    4.39,    4.39,    4.39,
  4.03,    4.03,    4.03,    4.03,
  4.23,    4.23,    4.23,    4.23,
  4.7,     4.7,     4.7,     4.7,
  4.36,    4.36,    4.36,    4.36,
  4.54,    4.54,    4.54,    4.54,
  4.58,    4.58,    4.58,    4.58,
  5.09,    5.09,    5.09,    5.09,
  5.35,    5.35,    5.35,    5.35,
  5,       5,       5,       5,
  5.71,    5.71,    5.71,    5.71,
  5.85,    5.85,    5.85,    5.85,
  6.24,    6.24,    6.24,    6.24,
  6.1,     6.1,     6.1,     6.1,
  6.31,    6.31,    6.31,    6.31,
  6.07,    6.07,    6.07,    6.07,
  4.92,    4.92,    4.92,    4.92,
  5.77,    5.77,    5.77,    5.77,
  5.03,    5.03,    5.03,    5.03,
  5.61,    5.61,    5.61,    5.61,
  4.69,    4.69,    4.69,    4.69,
  5.18,    5.18,    5.18,    5.18,
  5.24,    5.24,    5.24,    5.24,
  5.2,     5.2,     5.2,     5.2,
  5.45,    5.45,    5.45,    5.45,
  5.29,    5.29,    5.29,    5.29,
  5.51,    5.51,    5.51,    5.51,
  5.12,    5.12,    5.12,    5.12,
  5.55,    5.55,    5.55,    5.55,
  4.97,    4.97,    4.97,    4.97,
  5.07,    5.07,    5.07,    5.07,
  4.24,    4.24,    4.24,    4.24,
  4.62,    4.62,    4.62,    4.62,
  4.94,    4.94,    4.94,    4.94,
  5.1,     5.1,     5.1,     5.1,
  4.57,    4.57,    4.57,    4.57,
  5.56,    5.56,    5.56,    5.56,
  6.24,    6.24,    6.24,    6.24,
  5.44,    5.44,    5.44,    5.44,
  5.27,    5.27,    5.27,    5.27,
  5.26,    5.26,    5.26,    5.26,
  5.8,     5.8,     5.8,     5.8,
  5.77,    5.77,    5.77,    5.77,
  5.83,    5.83,    5.83,    5.83,
  5.09,    5.09,    5.09,    5.09,
  4.39,    4.39,    4.39,    4.39,
  3.93,    3.93,    3.93,    3.93,
  4.4,     4.4,     4.4,     4.4,
  3.86,    3.86,    3.86,    3.86,
  5.1,     5.1,     5.1,     5.1,
  5.51,    5.51,    5.51,    5.51,
  5.64,    5.64,    5.64,    5.64,
  5.64,    5.64,    5.64,    5.64,
  5.57,    5.57,    5.57,    5.57,
  4.71,    4.71,    4.71,    4.71,
  4.17,    4.17,    4.17,    4.17,
  4.43,    4.43,    4.43,    4.43,
  5.06,    5.06,    5.06,    5.06,
  5.55,    5.55,    5.55,    5.55,
  3.9,     3.9,     3.9,     3.9,
  4.03,    4.03,    4.03,    4.03,
  4.34,    4.34,    4.34,    4.34,
  5.25,    5.25,    5.25,    5.25,
  6.32,    6.32,    6.32,    6.32,
  6.15,    6.15,    6.15,    6.15,
  6.5,     6.5,     6.5,     6.5,
  7.1,     7.1,     7.1,     7.1,
  7.06,    7.06,    7.06,    7.06,
  6.5,     6.5,     6.5,     6.5,
  7.46,    7.46,    7.46,    7.46,
  6.69,    6.69,    6.69,    6.69,
  6.89,    6.89,    6.89,    6.89,
  6.74,    6.74,    6.74,    6.74,
  6.14,    6.14,    6.14,    6.14,
  6.7,     6.7,     6.7,     6.7,
  6.42,    6.42,    6.42,    6.42,
  6.23,    6.23,    6.23,    6.23,
  6.15,    6.15,    6.15,    6.15,
  6.71,    6.71,    6.71,    6.71,
  6.55,    6.55,    6.55,    6.55,
  6.55,    6.55,    6.55,    6.55,
  5.99,    5.99,    5.99,    5.99,
  5.21,    5.21,    5.21,    5.21,
  4.97,    4.97,    4.97,    4.97,
  4,       4,       4,       4,
  3.88,    3.88,    3.88,    3.88,
  3.54,    3.54,    3.54,    3.54,
  3.03,    3.03,    3.03,    3.03,
  3.34,    3.34,    3.34,    3.34,
  3.22,    3.22,    3.22,    3.22,
  3.1,     3.1,     3.1,     3.1,
  3.25,    3.25,    3.25,    3.25,
  2.93,    2.93,    2.93,    2.93,
  2.95,    2.95,    2.95,    2.95,
  2.52,    2.52,    2.52,    2.52,
  2.89,    2.89,    2.89,    2.89,
  3.05,    3.05,    3.05,    3.05,
  3.34,    3.34,    3.34,    3.34,
  3.47,    3.47,    3.47,    3.47,
  3.81,    3.81,    3.81,    3.81,
  4.64,    4.64,    4.64,    4.64,
  3.74,    3.74,    3.74,    3.74,
  3.46,    3.46,    3.46,    3.46,
  3.4,     3.4,     3.4,     3.4,
  4.39,    4.39,    4.39,    4.39,
  4.07,    4.07,    4.07,    4.07,
  3.95,    3.95,    3.95,    3.95,
  3.86,    3.86,    3.86,    3.86,
  3.96,    3.96,    3.96,    3.96,
  3.03,    3.03,    3.03,    3.03,
  4.08,    4.08,    4.08,    4.08,
  3.23,    3.23,    3.23,    3.23,
  2.45,    2.45,    2.45,    2.45,
  1.98,    1.98,    1.98,    1.98,
  1.98,    1.98,    1.98,    1.98,
  1.9,     1.9,     1.9,     1.9,
  1.7,     1.7,     1.7,     1.7,
  1.99,    1.99,    1.99,    1.99,
  2.52,    2.52,    2.52,    2.52,
  2.62,    2.62,    2.62,    2.62,
  1.96,    1.96,    1.96,    1.96,
  0.52,    0.52,    0.52,    0.52,
  1.61,    1.61,    1.61,    1.61,
  1.83,    1.83,    1.83,    1.83,
  2.13,    2.13,    2.13,    2.13,
  1.39,    1.39,    1.39,    1.39,
  1.63,    1.63,    1.63,    1.63,
  1.6,     1.6,     1.6,     1.6,
  1.9,     1.9,     1.9,     1.9,
  1.75,    1.75,    1.75,    1.75,
  2.2,     2.2,     2.2,     2.2,
  2.03,    2.03,    2.03,    2.03,
  2.14,    2.14,    2.14,    2.14,
  2.58,    2.58,    2.58,    2.58,
  2.07,    2.07,    2.07,    2.07,
  1.79,    1.79,    1.79,    1.79,
  2.41,    2.41,    2.41,    2.41,
  2.61,    2.61,    2.61,    2.61,
  2.6,     2.6,     2.6,     2.6,
  2.22,    2.22,    2.22,    2.22,
  2.17,    2.17,    2.17,    2.17,
  2.17,    2.17,    2.17,    2.17,
  2.16,    2.16,    2.16,    2.16,
  1.88,    1.88,    1.88,    1.88,
  1.81,    1.81,    1.81,    1.81,
  1.81,    1.81,    1.81,    1.81,
  2.38,    2.38,    2.38,    2.38,
  2.12,    2.12,    2.12,    2.12,
  2.79,    2.79,    2.79,    2.79,
  3.18,    3.18,    3.18,    3.18,
  3.62,    3.62,    3.62,    3.62,
  4.37,    4.37,    4.37,    4.37,
  3.63,    3.63,    3.63,    3.63,
  3.56,    3.56,    3.56,    3.56,
  4.11,    4.11,    4.11,    4.11,
  3.2,     3.2,     3.2,     3.2,
  3.59,    3.59,    3.59,    3.59,
  4.01,    4.01,    4.01,    4.01,
  3.05,    3.05,    3.05,    3.05,
  2.86,    2.86,    2.86,    2.86,
  2.79,    2.79,    2.79,    2.79,
  2.47,    2.47,    2.47,    2.47,
  2.2,     2.2,     2.2,     2.2,
  1.94,    1.94,    1.94,    1.94,
  1.94,    1.94,    1.94,    1.94,
  1.8,     1.8,     1.8,     1.8,
  1.75,    1.75,    1.75,    1.75,
  1.62,    1.62,    1.62,    1.62,
  1.5,     1.5,     1.5,     1.5,
  1.86,    1.86,    1.86,    1.86,
  1.81,    1.81,    1.81,    1.81,
  1.79,    1.79,    1.79,    1.79,
  1.41,    1.41,    1.41,    1.41,
  1.52,    1.52,    1.52,    1.52,
  1.32,    1.32,    1.32,    1.32,
  1.16,    1.16,    1.16,    1.16,
  1.77,    1.77,    1.77,    1.77,
  1.96,    1.96,    1.96,    1.96,
  1.91,    1.91,    1.91,    1.91,
  1.73,    1.73,    1.73,    1.73,
  1.91,    1.91,    1.91,    1.91,
  1.69,    1.69,    1.69,    1.69,
  1.53,    1.53,    1.53,    1.53,
  1.47,    1.47,    1.47,    1.47,
  1.38,    1.38,    1.38,    1.38,
  1.35,    1.35,    1.35,    1.35,
  1.56,    1.56,    1.56,    1.56,
  1.65,    1.65,    1.65,    1.65,
  1.45,    1.45,    1.45,    1.45,
  1.45,    1.45,    1.45,    1.45,
  1.59,    1.59,    1.59,    1.59,
  2.06,    2.06,    2.06,    2.06,
  2.06,    2.06,    2.06,    2.06,
  2.23,    2.23,    2.23,    2.23,
  2.12,    2.12,    2.12,    2.12,
  2.66,    2.66,    2.66,    2.66,
  2.37,    2.37,    2.37,    2.37,
  3.41,    3.41,    3.41,    3.41,
  2.61,    2.61,    2.61,    2.61,
  3.57,    3.57,    3.57,    3.57,
  3.29,    3.29,    3.29,    3.29,
  3.44,    3.44,    3.44,    3.44,
  3.61,    3.61,    3.61,    3.61,
  3.44,    3.44,    3.44,    3.44,
  3.62,    3.62,    3.62,    3.62,
  3.24,    3.24,    3.24,    3.24,
  2.86,    2.86,    2.86,    2.86,
  2.83,    2.83,    2.83,    2.83,
  3.08,    3.08,    3.08,    3.08,
  2.77,    2.77,    2.77,    2.77,
  2.86,    2.86,    2.86,    2.86,
  2.83,    2.83,    2.83,    2.83,
  3.55,    3.55,    3.55,    3.55,
  3.49,    3.49,    3.49,    3.49,
  3.36,    3.36,    3.36,    3.36,
  3.08,    3.08,    3.08,    3.08,
  3.06,    3.06,    3.06,    3.06,
  3.16,    3.16,    3.16,    3.16,
  3.66,    3.66,    3.66,    3.66,
  3.43,    3.43,    3.43,    3.43,
  3.67,    3.67,    3.67,    3.67,
  3.89,    3.89,    3.89,    3.89,
  3.91,    3.91,    3.91,    3.91,
  3.48,    3.48,    3.48,    3.48,
  3.79,    3.79,    3.79,    3.79,
  3.94,    3.94,    3.94,    3.94,
  3.89,    3.89,    3.89,    3.89,
  3.85,    3.85,    3.85,    3.85,
  2.85,    2.85,    2.85,    2.85,
  3.16,    3.16,    3.16,    3.16,
  3.38,    3.38,    3.38,    3.38,
  3.01,    3.01,    3.01,    3.01,
  2.94,    2.94,    2.94,    2.94,
  2.86,    2.86,    2.86,    2.86,
  3,       3,       3,       3,
  2.57,    2.57,    2.57,    2.57,
  2.7,     2.7,     2.7,     2.7,
  2.61,    2.61,    2.61,    2.61,
  2.92,    2.92,    2.92,    2.92,
  2.91,    2.91,    2.91,    2.91,
  2.73,    2.73,    2.73,    2.73,
  2.54,    2.54,    2.54,    2.54,
  2.77,    2.77,    2.77,    2.77,
  2.99,    2.99,    2.99,    2.99,
  2.78,    2.78,    2.78,    2.78,
  3.59,    3.59,    3.59,    3.59,
  3.26,    3.26,    3.26,    3.26,
  3.49,    3.49,    3.49,    3.49,
  3.63,    3.63,    3.63,    3.63,
  3.56,    3.56,    3.56,    3.56,
  4.17,    4.17,    4.17,    4.17,
  4.09,    4.09,    4.09,    4.09,
  4.18,    4.18,    4.18,    4.18,
  2.95,    2.95,    2.95,    2.95,
  3.23,    3.23,    3.23,    3.23,
  3.24,    3.24,    3.24,    3.24,
  3.32,    3.32,    3.32,    3.32,
  3.51,    3.51,    3.51,    3.51,
  3.29,    3.29,    3.29,    3.29,
  3.54,    3.54,    3.54,    3.54,
  3.72,    3.72,    3.72,    3.72,
  4.29,    4.29,    4.29,    4.29,
  4.41,    4.41,    4.41,    4.41,
  4.46,    4.46,    4.46,    4.46,
  4.4,     4.4,     4.4,     4.4,
  4.27,    4.27,    4.27,    4.27,
  4.38,    4.38,    4.38,    4.38,
  4.57,    4.57,    4.57,    4.57,
  5.01,    5.01,    5.01,    5.01,
  5.22,    5.22,    5.22,    5.22,
  5.24,    5.24,    5.24,    5.24,
  4.51,    4.51,    4.51,    4.51,
  4.83,    4.83,    4.83,    4.83,
  4.72,    4.72,    4.72,    4.72,
  5,       5,       5,       5,
  5.03,    5.03,    5.03,    5.03,
  5.02,    5.02,    5.02,    5.02,
  4.96,    4.96,    4.96,    4.96,
  5.42,    5.42,    5.42,    5.42,
  5.21,    5.21,    5.21,    5.21,
  4.97,    4.97,    4.97,    4.97,
  4.82,    4.82,    4.82,    4.82,
  5.3,     5.3,     5.3,     5.3,
  4.57,    4.57,    4.57,    4.57,
  4.71,    4.71,    4.71,    4.71,
  4.78,    4.78,    4.78,    4.78,
  4.38,    4.38,    4.38,    4.38,
  4.15,    4.15,    4.15,    4.15,
  4.35,    4.35,    4.35,    4.35,
  5.1,     5.1,     5.1,     5.1,
  6.34,    6.34,    6.34,    6.34,
  6.3,     6.3,     6.3,     6.3,
  5.64,    5.64,    5.64,    5.64,
  6.07,    6.07,    6.07,    6.07,
  6.53,    6.53,    6.53,    6.53,
  8.79,    8.79,    8.79,    8.79,
  7.41,    7.41,    7.41,    7.41,
  7.64,    7.64,    7.64,    7.64,
  7.06,    7.06,    7.06,    7.06,
  7.41,    7.41,    7.41,    7.41,
  7.76,    7.76,    7.76,    7.76,
  7.87,    7.87,    7.87,    7.87,
  6.82,    6.82,    6.82,    6.82,
  5.47,    5.47,    5.47,    5.47,
  5.52,    5.52,    5.52,    5.52,
  4.49,    4.49,    4.49,    4.49,
  3.88,    3.88,    3.88,    3.88,
  2.83,    2.83,    2.83,    2.83,
  2.54,    2.54,    2.54,    2.54,
  2.76,    2.76,    2.76,    2.76,
  3.35,    3.35,    3.35,    3.35,
  4.54,    4.54,    4.54,    4.54,
  4.61,    4.61,    4.61,    4.61,
  5.72,    5.72,    5.72,    5.72,
  5.47,    5.47,    5.47,    5.47,
  5.44,    5.44,    5.44,    5.44,
  4.92,    4.92,    4.92,    4.92,
  4.87,    4.87,    4.87,    4.87,
  4.84,    4.84,    4.84,    4.84,
  4.99,    4.99,    4.99,    4.99,
  4.81,    4.81,    4.81,    4.81,
  4.6,     4.6,     4.6,     4.6,
  4.44,    4.44,    4.44,    4.44,
  5,       5,       5,       5,
  4.2,     4.2,     4.2,     4.2,
  4.67,    4.67,    4.67,    4.67,
  4.8,     4.8,     4.8,     4.8,
  4,       4,       4,       4,
  4.1,     4.1,     4.1,     4.1,
  3.59,    3.59,    3.59,    3.59,
  2.64,    2.64,    2.64,    2.64,
  2.46,    2.46,    2.46,    2.46,
  2.32,    2.32,    2.32,    2.32,
  2.77,    2.77,    2.77,    2.77,
  3.06,    3.06,    3.06,    3.06,
  2.65,    2.65,    2.65,    2.65,
  2.56,    2.56,    2.56,    2.56,
  2.9,     2.9,     2.9,     2.9,
  3.27,    3.27,    3.27,    3.27,
  3.53,    3.53,    3.53,    3.53,
  3.8,     3.8,     3.8,     3.8,
  3.88,    3.88,    3.88,    3.88,
  4.41,    4.41,    4.41,    4.41,
  4.4,     4.4,     4.4,     4.4,
  4.14,    4.14,    4.14,    4.14,
  4.3,     4.3,     4.3,     4.3,
  4.76,    4.76,    4.76,    4.76,
  4.49,    4.49,    4.49,    4.49,
  4.64,    4.64,    4.64,    4.64,
  5.05,    5.05,    5.05,    5.05,
  4.82,    4.82,    4.82,    4.82,
  5.48,    5.48,    5.48,    5.48,
  5.69,    5.69,    5.69,    5.69,
  5.72,    5.72,    5.72,    5.72,
  6.08,    6.08,    6.08,    6.08,
  6.24,    6.24,    6.24,    6.24,
  6.26,    6.26,    6.26,    6.26,
  6.24,    6.24,    6.24,    6.24,
  6.25,    6.25,    6.25,    6.25,
  6.24,    6.24,    6.24,    6.24,
  6.77,    6.77,    6.77,    6.77,
  6.89,    6.89,    6.89,    6.89,
  6.65,    6.65,    6.65,    6.65,
  6.42,    6.42,    6.42,    6.42,
  6.8,     6.8,     6.8,     6.8,
  6.54,    6.54,    6.54,    6.54,
  7.89,    7.89,    7.89,    7.89,
  7.7,     7.7,     7.7,     7.7,
  7.81,    7.81,    7.81,    7.81,
  8.54,    8.54,    8.54,    8.54,
  8.7,     8.7,     8.7,     8.7,
  6.63,    6.63,    6.63,    6.63,
  7.59,    7.59,    7.59,    7.59,
  7.98,    7.98,    7.98,    7.98,
  7.35,    7.35,    7.35,    7.35,
  6.59,    6.59,    6.59,    6.59,
  6.64,    6.64,    6.64,    6.64,
  5.89,    5.89,    5.89,    5.89,
  6.02,    6.02,    6.02,    6.02,
  6.05,    6.05,    6.05,    6.05,
  6.03,    6.03,    6.03,    6.03,
  6.32,    6.32,    6.32,    6.32,
  5.82,    5.82,    5.82,    5.82,
  5.27,    5.27,    5.27,    5.27,
  5.57,    5.57,    5.57,    5.57,
  4.91,    4.91,    4.91,    4.91,
  6.19,    6.19,    6.19,    6.19,
  6.17,    6.17,    6.17,    6.17,
  5.64,    5.64,    5.64,    5.64,
  5.81,    5.81,    5.81,    5.81,
  4.34,    4.34,    4.34,    4.34,
  4.77,    4.77,    4.77,    4.77,
  5.56,    5.56,    5.56,    5.56,
  5.63,    5.63,    5.63,    5.63,
  5.96,    5.96,    5.96,    5.96,
  5.71,    5.71,    5.71,    5.71,
  6.02,    6.02,    6.02,    6.02,
  5.41,    5.41,    5.41,    5.41,
  5.6,     5.6,     5.6,     5.6,
  6.28,    6.28,    6.28,    6.28,
  5.25,    5.25,    5.25,    5.25,
  5.49,    5.49,    5.49,    5.49,
  4.79,    4.79,    4.79,    4.79,
  5.23,    5.23,    5.23,    5.23,
  4.94,    4.94,    4.94,    4.94,
  5.56,    5.56,    5.56,    5.56,
  5.61,    5.61,    5.61,    5.61,
  5.79,    5.79,    5.79,    5.79,
  6.53,    6.53,    6.53,    6.53,
  6.63,    6.63,    6.63,    6.63,
  5.32,    5.32,    5.32,    5.32,
  5.42,    5.42,    5.42,    5.42,
  6.03,    6.03,    6.03,    6.03,
  6.15,    6.15,    6.15,    6.15,
  5.35,    5.35,    5.35,    5.35,
  6.03,    6.03,    6.03,    6.03,
  7.06,    7.06,    7.06,    7.06,
  6.65,    6.65,    6.65,    6.65,
  6.18,    6.18,    6.18,    6.18,
  5.9,     5.9,     5.9,     5.9,
  5.72,    5.72,    5.72,    5.72,
  5.93,    5.93,    5.93,    5.93,
  5.74,    5.74,    5.74,    5.74,
  5.59,    5.59,    5.59,    5.59,
  5.55,    5.55,    5.55,    5.55,
  5.73,    5.73,    5.73,    5.73,
  7.17,    7.17,    7.17,    7.17,
  6.56,    6.56,    6.56,    6.56,
  6.46,    6.46,    6.46,    6.46,
  6.17,    6.17,    6.17,    6.17,
  6.21,    6.21,    6.21,    6.21,
  6.81,    6.81,    6.81,    6.81,
  6.19,    6.19,    6.19,    6.19,
  6.82,    6.82,    6.82,    6.82,
  6.37,    6.37,    6.37,    6.37,
  6.71,    6.71,    6.71,    6.71,
  6.21,    6.21,    6.21,    6.21,
  6.06,    6.06,    6.06,    6.06,
  5.68,    5.68,    5.68,    5.68,
  5.37,    5.37,    5.37,    5.37,
  5.44,    5.44,    5.44,    5.44,
  5.83,    5.83,    5.83,    5.83,
  5.43,    5.43,    5.43,    5.43,
  4.7,     4.7,     4.7,     4.7,
  5.31,    5.31,    5.31,    5.31,
  4.8,     4.8,     4.8,     4.8,
  5.11,    5.11,    5.11,    5.11,
  4.1,     4.1,     4.1,     4.1,
  4.52,    4.52,    4.52,    4.52,
  4.58,    4.58,    4.58,    4.58,
  3.36,    3.36,    3.36,    3.36,
  2.52,    2.52,    2.52,    2.52,
  2.76,    2.76,    2.76,    2.76,
  3.07,    3.07,    3.07,    3.07,
  2.36,    2.36,    2.36,    2.36,
  2.57,    2.57,    2.57,    2.57,
  2.19,    2.19,    2.19,    2.19,
  2.61,    2.61,    2.61,    2.61,
  2.55,    2.55,    2.55,    2.55,
  2.43,    2.43,    2.43,    2.43,
  2.54,    2.54,    2.54,    2.54,
  2.46,    2.46,    2.46,    2.46,
  2.84,    2.84,    2.84,    2.84,
  2.6,     2.6,     2.6,     2.6,
  2.72,    2.72,    2.72,    2.72,
  2.7,     2.7,     2.7,     2.7,
  2.41,    2.41,    2.41,    2.41,
  2.48,    2.48,    2.48,    2.48,
  2.35,    2.35,    2.35,    2.35,
  3.15,    3.15,    3.15,    3.15,
  3.49,    3.49,    3.49,    3.49,
  3.32,    3.32,    3.32,    3.32,
  3.07,    3.07,    3.07,    3.07,
  3.23,    3.23,    3.23,    3.23,
  3.21,    3.21,    3.21,    3.21,
  3.21,    3.21,    3.21,    3.21,
  3.66,    3.66,    3.66,    3.66,
  3.44,    3.44,    3.44,    3.44,
  3.59,    3.59,    3.59,    3.59,
  3.57,    3.57,    3.57,    3.57,
  3.76,    3.76,    3.76,    3.76,
  3.29,    3.29,    3.29,    3.29,
  3.28,    3.28,    3.28,    3.28,
  3.35,    3.35,    3.35,    3.35,
  3.18,    3.18,    3.18,    3.18,
  3.44,    3.44,    3.44,    3.44,
  3.26,    3.26,    3.26,    3.26,
  3.49,    3.49,    3.49,    3.49,
  3.18,    3.18,    3.18,    3.18,
  3.43,    3.43,    3.43,    3.43,
  3.32,    3.32,    3.32,    3.32,
  3.81,    3.81,    3.81,    3.81,
  3.66,    3.66,    3.66,    3.66,
  3.2,     3.2,     3.2,     3.2,
  3.32,    3.32,    3.32,    3.32,
  3.28,    3.28,    3.28,    3.28,
  2.94,    2.94,    2.94,    2.94,
  2.84,    2.84,    2.84,    2.84,
  2.46,    2.46,    2.46,    2.46,
  2.16,    2.16,    2.16,    2.16,
  2.03,    2.03,    2.03,    2.03,
  1.87,    1.87,    1.87,    1.87,
  1.53,    1.53,    1.53,    1.53,
  2.51,    2.51,    2.51,    2.51,
  3.08,    3.08,    3.08,    3.08,
  2.67,    2.67,    2.67,    2.67,
  2.9,     2.9,     2.9,     2.9,
  2.64,    2.64,    2.64,    2.64,
  2.78,    2.78,    2.78,    2.78,
  3.38,    3.38,    3.38,    3.38,
  3.09,    3.09,    3.09,    3.09,
  2.92,    2.92,    2.92,    2.92,
  2.96,    2.96,    2.96,    2.96,
  2.93,    2.93,    2.93,    2.93,
  2.66,    2.66,    2.66,    2.66,
  2.63,    2.63,    2.63,    2.63,
  2.28,    2.28,    2.28,    2.28,
  2.36,    2.36,    2.36,    2.36,
  2.71,    2.71,    2.71,    2.71,
  2.78,    2.78,    2.78,    2.78,
  2.87,    2.87,    2.87,    2.87,
  2.54,    2.54,    2.54,    2.54,
  2.34,    2.34,    2.34,    2.34,
  1.97,    1.97,    1.97,    1.97,
  2.2,     2.2,     2.2,     2.2,
  2.65,    2.65,    2.65,    2.65,
  3.37,    3.37,    3.37,    3.37,
  3.12,    3.12,    3.12,    3.12,
  3.26,    3.26,    3.26,    3.26,
  3.56,    3.56,    3.56,    3.56,
  3.4,     3.4,     3.4,     3.4,
  3.42,    3.42,    3.42,    3.42,
  3.64,    3.64,    3.64,    3.64,
  3.86,    3.86,    3.86,    3.86,
  4.09,    4.09,    4.09,    4.09,
  4.32,    4.32,    4.32,    4.32,
  4.47,    4.47,    4.47,    4.47,
  5.08,    5.08,    5.08,    5.08,
  4.46,    4.46,    4.46,    4.46,
  5.05,    5.05,    5.05,    5.05,
  4.92,    4.92,    4.92,    4.92,
  4.26,    4.26,    4.26,    4.26,
  4.27,    4.27,    4.27,    4.27,
  3.94,    3.94,    3.94,    3.94,
  4.03,    4.03,    4.03,    4.03,
  4.07,    4.07,    4.07,    4.07,
  3.78,    3.78,    3.78,    3.78,
  4.09,    4.09,    4.09,    4.09,
  4.5,     4.5,     4.5,     4.5,
  4.51,    4.51,    4.51,    4.51,
  4.53,    4.53,    4.53,    4.53,
  4.52,    4.52,    4.52,    4.52,
  3.63,    3.63,    3.63,    3.63,
  4.14,    4.14,    4.14,    4.14,
  3.94,    3.94,    3.94,    3.94,
  4,       4,       4,       4,
  4.5,     4.5,     4.5,     4.5,
  4.88,    4.88,    4.88,    4.88,
  5.44,    5.44,    5.44,    5.44,
  5.12,    5.12,    5.12,    5.12,
  5.07,    5.07,    5.07,    5.07,
  5.42,    5.42,    5.42,    5.42,
  6.12,    6.12,    6.12,    6.12,
  5.41,    5.41,    5.41,    5.41,
  5.76,    5.76,    5.76,    5.76,
  5.41,    5.41,    5.41,    5.41,
  5.37,    5.37,    5.37,    5.37,
  5.52,    5.52,    5.52,    5.52,
  5.99,    5.99,    5.99,    5.99,
  5.92,    5.92,    5.92,    5.92,
  5.73,    5.73,    5.73,    5.73,
  5.64,    5.64,    5.64,    5.64,
  5.18,    5.18,    5.18,    5.18,
  5.4,     5.4,     5.4,     5.4,
  5.55,    5.55,    5.55,    5.55,
  5.3,     5.3,     5.3,     5.3,
  4.76,    4.76,    4.76,    4.76,
  3.62,    3.62,    3.62,    3.62,
  3.35,    3.35,    3.35,    3.35,
  4.82,    4.82,    4.82,    4.82,
  4.31,    4.31,    4.31,    4.31,
  3.3,     3.3,     3.3,     3.3,
  3.5,     3.5,     3.5,     3.5,
  4.2,     4.2,     4.2,     4.2,
  3.63,    3.63,    3.63,    3.63,
  3.95,    3.95,    3.95,    3.95,
  4.89,    4.89,    4.89,    4.89,
  4.47,    4.47,    4.47,    4.47,
  3.64,    3.64,    3.64,    3.64,
  4.13,    4.13,    4.13,    4.13,
  3.94,    3.94,    3.94,    3.94,
  4.54,    4.54,    4.54,    4.54,
  4.17,    4.17,    4.17,    4.17,
  4.34,    4.34,    4.34,    4.34,
  4.19,    4.19,    4.19,    4.19,
  4.39,    4.39,    4.39,    4.39,
  4.39,    4.39,    4.39,    4.39,
  4.71,    4.71,    4.71,    4.71,
  5.23,    5.23,    5.23,    5.23,
  5.21,    5.21,    5.21,    5.21,
  4.65,    4.65,    4.65,    4.65,
  4.62,    4.62,    4.62,    4.62,
  4.8,     4.8,     4.8,     4.8,
  6.55,    6.55,    6.55,    6.55,
  6.94,    6.94,    6.94,    6.94,
  7.69,    7.69,    7.69,    7.69,
  7.91,    7.91,    7.91,    7.91,
  8.3,     8.3,     8.3,     8.3,
  8.1,     8.1,     8.1,     8.1,
  8.6,     8.6,     8.6,     8.6,
  6.82,    6.82,    6.82,    6.82,
  8.56,    8.56,    8.56,    8.56,
  8.65,    8.65,    8.65,    8.65,
  9.66,    9.66,    9.66,    9.66,
  9.37,    9.37,    9.37,    9.37,
  8.7,     8.7,     8.7,     8.7,
  7.65,    7.65,    7.65,    7.65,
  6.48,    6.48,    6.48,    6.48,
  8.19,    8.19,    8.19,    8.19,
  7.58,    7.58,    7.58,    7.58,
  7.13,    7.13,    7.13,    7.13,
  5.85,    5.85,    5.85,    5.85,
  6.04,    6.04,    6.04,    6.04,
  7.2,     7.2,     7.2,     7.2,
  7.36,    7.36,    7.36,    7.36,
  8.1,     8.1,     8.1,     8.1,
  7.41,    7.41,    7.41,    7.41,
  7.03,    7.03,    7.03,    7.03,
  6.88,    6.88,    6.88,    6.88,
  8.01,    8.01,    8.01,    8.01,
  7.86,    7.86,    7.86,    7.86,
  7.99,    7.99,    7.99,    7.99,
  7.64,    7.64,    7.64,    7.64,
  7.08,    7.08,    7.08,    7.08,
  8.16,    8.16,    8.16,    8.16,
  7.56,    7.56,    7.56,    7.56,
  8.1,     8.1,     8.1,     8.1,
  7.99,    7.99,    7.99,    7.99,
  7.84,    7.84,    7.84,    7.84,
  7.44,    7.44,    7.44,    7.44,
  6.94,    6.94,    6.94,    6.94,
  7.74,    7.74,    7.74,    7.74,
  6.73,    6.73,    6.73,    6.73,
  6.53,    6.53,    6.53,    6.53,
  6.66,    6.66,    6.66,    6.66,
  5.86,    5.86,    5.86,    5.86,
  5.75,    5.75,    5.75,    5.75,
  5.12,    5.12,    5.12,    5.12,
  5.43,    5.43,    5.43,    5.43,
  5.55,    5.55,    5.55,    5.55,
  4.99,    4.99,    4.99,    4.99,
  4.4,     4.4,     4.4,     4.4,
  5.36,    5.36,    5.36,    5.36,
  4.22,    4.22,    4.22,    4.22,
  5.43,    5.43,    5.43,    5.43,
  5.41,    5.41,    5.41,    5.41,
  4.97,    4.97,    4.97,    4.97,
  5.44,    5.44,    5.44,    5.44,
  5.54,    5.54,    5.54,    5.54,
  5.61,    5.61,    5.61,    5.61,
  5.22,    5.22,    5.22,    5.22,
  5.86,    5.86,    5.86,    5.86,
  5.02,    5.02,    5.02,    5.02,
  5.48,    5.48,    5.48,    5.48,
  5.43,    5.43,    5.43,    5.43,
  5.01,    5.01,    5.01,    5.01,
  5.18,    5.18,    5.18,    5.18,
  5.21,    5.21,    5.21,    5.21,
  4.85,    4.85,    4.85,    4.85,
  5.23,    5.23,    5.23,    5.23,
  5.28,    5.28,    5.28,    5.28,
  5.07,    5.07,    5.07,    5.07,
  4.5,     4.5,     4.5,     4.5,
  5.91,    5.91,    5.91,    5.91,
  4.86,    4.86,    4.86,    4.86,
  5.32,    5.32,    5.32,    5.32,
  5.61,    5.61,    5.61,    5.61,
  4.67,    4.67,    4.67,    4.67,
  5.05,    5.05,    5.05,    5.05,
  5.91,    5.91,    5.91,    5.91,
  5.28,    5.28,    5.28,    5.28,
  4.04,    4.04,    4.04,    4.04,
  6.2,     6.2,     6.2,     6.2,
  6.79,    6.79,    6.79,    6.79,
  6.15,    6.15,    6.15,    6.15,
  5.65,    5.65,    5.65,    5.65,
  4.89,    4.89,    4.89,    4.89,
  3.57,    3.57,    3.57,    3.57,
  3.9,     3.9,     3.9,     3.9,
  4.71,    4.71,    4.71,    4.71,
  3.94,    3.94,    3.94,    3.94,
  3.77,    3.77,    3.77,    3.77,
  3.87,    3.87,    3.87,    3.87,
  4.78,    4.78,    4.78,    4.78,
  4.1,     4.1,     4.1,     4.1,
  3.85,    3.85,    3.85,    3.85,
  3.81,    3.81,    3.81,    3.81,
  3.69,    3.69,    3.69,    3.69,
  3.82,    3.82,    3.82,    3.82,
  4.21,    4.21,    4.21,    4.21,
  4.18,    4.18,    4.18,    4.18,
  4.03,    4.03,    4.03,    4.03,
  3.7,     3.7,     3.7,     3.7,
  3.73,    3.73,    3.73,    3.73,
  3.68,    3.68,    3.68,    3.68,
  4.19,    4.19,    4.19,    4.19,
  4.53,    4.53,    4.53,    4.53,
  4.69,    4.69,    4.69,    4.69,
  3.49,    3.49,    3.49,    3.49,
  3.37,    3.37,    3.37,    3.37,
  2.78,    2.78,    2.78,    2.78,
  2.68,    2.68,    2.68,    2.68,
  2.1,     2.1,     2.1,     2.1,
  1.95,    1.95,    1.95,    1.95,
  2.08,    2.08,    2.08,    2.08,
  2.41,    2.41,    2.41,    2.41,
  2.2,     2.2,     2.2,     2.2,
  2.16,    2.16,    2.16,    2.16,
  1.88,    1.88,    1.88,    1.88,
  1.92,    1.92,    1.92,    1.92,
  1.68,    1.68,    1.68,    1.68,
  2.23,    2.23,    2.23,    2.23,
  1.96,    1.96,    1.96,    1.96,
  2.19,    2.19,    2.19,    2.19,
  2.23,    2.23,    2.23,    2.23,
  2.4,     2.4,     2.4,     2.4,
  2.92,    2.92,    2.92,    2.92,
  2.69,    2.69,    2.69,    2.69,
  2.98,    2.98,    2.98,    2.98,
  2.73,    2.73,    2.73,    2.73,
  3.28,    3.28,    3.28,    3.28,
  3.63,    3.63,    3.63,    3.63,
  3.31,    3.31,    3.31,    3.31,
  4.18,    4.18,    4.18,    4.18,
  3.53,    3.53,    3.53,    3.53,
  2.85,    2.85,    2.85,    2.85,
  2.74,    2.74,    2.74,    2.74,
  2.54,    2.54,    2.54,    2.54,
  2.85,    2.85,    2.85,    2.85,
  2.31,    2.31,    2.31,    2.31,
  2.38,    2.38,    2.38,    2.38,
  2.03,    2.03,    2.03,    2.03,
  2.04,    2.04,    2.04,    2.04,
  2.08,    2.08,    2.08,    2.08,
  2.66,    2.66,    2.66,    2.66,
  3.6,     3.6,     3.6,     3.6,
  3.73,    3.73,    3.73,    3.73,
  3.66,    3.66,    3.66,    3.66,
  3.44,    3.44,    3.44,    3.44,
  3.54,    3.54,    3.54,    3.54,
  3.57,    3.57,    3.57,    3.57,
  3.65,    3.65,    3.65,    3.65,
  3.53,    3.53,    3.53,    3.53,
  3.31,    3.31,    3.31,    3.31,
  3.41,    3.41,    3.41,    3.41,
  3.37,    3.37,    3.37,    3.37,
  3.51,    3.51,    3.51,    3.51,
  4.1,     4.1,     4.1,     4.1,
  4.03,    4.03,    4.03,    4.03,
  4.4,     4.4,     4.4,     4.4,
  4.03,    4.03,    4.03,    4.03,
  3.73,    3.73,    3.73,    3.73,
  3.85,    3.85,    3.85,    3.85,
  3.62,    3.62,    3.62,    3.62,
  3.65,    3.65,    3.65,    3.65,
  3.76,    3.76,    3.76,    3.76,
  3.88,    3.88,    3.88,    3.88,
  4.01,    4.01,    4.01,    4.01,
  5.07,    5.07,    5.07,    5.07,
  5.2,     5.2,     5.2,     5.2,
  4.48,    4.48,    4.48,    4.48,
  4.8,     4.8,     4.8,     4.8,
  4.96,    4.96,    4.96,    4.96,
  4.56,    4.56,    4.56,    4.56,
  3.79,    3.79,    3.79,    3.79,
  4.27,    4.27,    4.27,    4.27,
  4.73,    4.73,    4.73,    4.73,
  4.18,    4.18,    4.18,    4.18,
  4.03,    4.03,    4.03,    4.03,
  3.79,    3.79,    3.79,    3.79,
  4.23,    4.23,    4.23,    4.23,
  3.7,     3.7,     3.7,     3.7,
  3.2,     3.2,     3.2,     3.2,
  3.72,    3.72,    3.72,    3.72,
  3.81,    3.81,    3.81,    3.81,
  3,       3,       3,       3,
  2.32,    2.32,    2.32,    2.32,
  2.78,    2.78,    2.78,    2.78,
  2.92,    2.92,    2.92,    2.92,
  2.98,    2.98,    2.98,    2.98,
  3.04,    3.04,    3.04,    3.04,
  3.13,    3.13,    3.13,    3.13,
  3.05,    3.05,    3.05,    3.05,
  2.68,    2.68,    2.68,    2.68,
  3.18,    3.18,    3.18,    3.18,
  3.19,    3.19,    3.19,    3.19,
  2.83,    2.83,    2.83,    2.83,
  2.49,    2.49,    2.49,    2.49,
  2.2,     2.2,     2.2,     2.2,
  2.31,    2.31,    2.31,    2.31,
  2.61,    2.61,    2.61,    2.61,
  2.55,    2.55,    2.55,    2.55,
  2.91,    2.91,    2.91,    2.91,
  2.84,    2.84,    2.84,    2.84,
  2.51,    2.51,    2.51,    2.51,
  2.55,    2.55,    2.55,    2.55,
  1.92,    1.92,    1.92,    1.92,
  2.08,    2.08,    2.08,    2.08,
  2.05,    2.05,    2.05,    2.05,
  2.06,    2.06,    2.06,    2.06,
  2,       2,       2,       2,
  2.11,    2.11,    2.11,    2.11,
  2.04,    2.04,    2.04,    2.04,
  2.07,    2.07,    2.07,    2.07,
  2.31,    2.31,    2.31,    2.31,
  2.22,    2.22,    2.22,    2.22,
  2.38,    2.38,    2.38,    2.38,
  2.75,    2.75,    2.75,    2.75,
  2.99,    2.99,    2.99,    2.99,
  2.92,    2.92,    2.92,    2.92,
  3.4,     3.4,     3.4,     3.4,
  3.87,    3.87,    3.87,    3.87,
  3.78,    3.78,    3.78,    3.78,
  3.6,     3.6,     3.6,     3.6,
  4.25,    4.25,    4.25,    4.25,
  4.02,    4.02,    4.02,    4.02,
  3.36,    3.36,    3.36,    3.36,
  4.17,    4.17,    4.17,    4.17,
  4.69,    4.69,    4.69,    4.69,
  5.23,    5.23,    5.23,    5.23,
  5.05,    5.05,    5.05,    5.05,
  4.46,    4.46,    4.46,    4.46,
  4.23,    4.23,    4.23,    4.23,
  3.08,    3.08,    3.08,    3.08,
  2.4,     2.4,     2.4,     2.4,
  2.55,    2.55,    2.55,    2.55,
  3.04,    3.04,    3.04,    3.04,
  3.41,    3.41,    3.41,    3.41,
  3.31,    3.31,    3.31,    3.31,
  3.65,    3.65,    3.65,    3.65,
  4.5,     4.5,     4.5,     4.5,
  4.54,    4.54,    4.54,    4.54,
  4.21,    4.21,    4.21,    4.21,
  4.2,     4.2,     4.2,     4.2,
  4.28,    4.28,    4.28,    4.28,
  4.78,    4.78,    4.78,    4.78,
  4.69,    4.69,    4.69,    4.69,
  4.41,    4.41,    4.41,    4.41,
  4.35,    4.35,    4.35,    4.35,
  4.62,    4.62,    4.62,    4.62,
  4.61,    4.61,    4.61,    4.61,
  4.2,     4.2,     4.2,     4.2,
  4.51,    4.51,    4.51,    4.51,
  4.93,    4.93,    4.93,    4.93,
  4.78,    4.78,    4.78,    4.78,
  4.31,    4.31,    4.31,    4.31,
  4.31,    4.31,    4.31,    4.31,
  4.13,    4.13,    4.13,    4.13,
  4.27,    4.27,    4.27,    4.27,
  4.54,    4.54,    4.54,    4.54,
  5.34,    5.34,    5.34,    5.34,
  4.95,    4.95,    4.95,    4.95,
  5.22,    5.22,    5.22,    5.22,
  4.81,    4.81,    4.81,    4.81,
  4.86,    4.86,    4.86,    4.86,
  5.05,    5.05,    5.05,    5.05,
  5.92,    5.92,    5.92,    5.92,
  5.85,    5.85,    5.85,    5.85,
  6.85,    6.85,    6.85,    6.85,
  6.69,    6.69,    6.69,    6.69,
  6.07,    6.07,    6.07,    6.07,
  5.59,    5.59,    5.59,    5.59,
  5.1,     5.1,     5.1,     5.1,
  5.28,    5.28,    5.28,    5.28,
  4.84,    4.84,    4.84,    4.84,
  5.51,    5.51,    5.51,    5.51,
  5.04,    5.04,    5.04,    5.04,
  5.31,    5.31,    5.31,    5.31,
  3.95,    3.95,    3.95,    3.95,
  3.26,    3.26,    3.26,    3.26,
  2.95,    2.95,    2.95,    2.95,
  2.5,     2.5,     2.5,     2.5,
  2.53,    2.53,    2.53,    2.53,
  2.49,    2.49,    2.49,    2.49,
  2.44,    2.44,    2.44,    2.44,
  2.72,    2.72,    2.72,    2.72,
  2.67,    2.67,    2.67,    2.67,
  2.62,    2.62,    2.62,    2.62,
  2.45,    2.45,    2.45,    2.45,
  2.64,    2.64,    2.64,    2.64,
  2.58,    2.58,    2.58,    2.58,
  2.64,    2.64,    2.64,    2.64,
  2.73,    2.73,    2.73,    2.73,
  2.61,    2.61,    2.61,    2.61,
  2.46,    2.46,    2.46,    2.46,
  2.25,    2.25,    2.25,    2.25,
  2.56,    2.56,    2.56,    2.56,
  2.04,    2.04,    2.04,    2.04,
  1.94,    1.94,    1.94,    1.94,
  2.03,    2.03,    2.03,    2.03,
  1.97,    1.97,    1.97,    1.97,
  2.02,    2.02,    2.02,    2.02,
  2.19,    2.19,    2.19,    2.19,
  2.26,    2.26,    2.26,    2.26,
  2.47,    2.47,    2.47,    2.47,
  2.57,    2.57,    2.57,    2.57,
  2.57,    2.57,    2.57,    2.57,
  2.4,     2.4,     2.4,     2.4,
  2.4,     2.4,     2.4,     2.4,
  2.24,    2.24,    2.24,    2.24,
  2.67,    2.67,    2.67,    2.67,
  2.25,    2.25,    2.25,    2.25,
  2.05,    2.05,    2.05,    2.05,
  1.75,    1.75,    1.75,    1.75,
  2.42,    2.42,    2.42,    2.42,
  2.34,    2.34,    2.34,    2.34,
  2.44,    2.44,    2.44,    2.44,
  2.62,    2.62,    2.62,    2.62,
  2.93,    2.93,    2.93,    2.93,
  2.47,    2.47,    2.47,    2.47,
  2.82,    2.82,    2.82,    2.82,
  3.08,    3.08,    3.08,    3.08,
  2.94,    2.94,    2.94,    2.94,
  2.75,    2.75,    2.75,    2.75,
  2.52,    2.52,    2.52,    2.52,
  2.42,    2.42,    2.42,    2.42,
  1.57,    1.57,    1.57,    1.57,
  1.17,    1.17,    1.17,    1.17,
  1.35,    1.35,    1.35,    1.35,
  1.32,    1.32,    1.32,    1.32,
  1.69,    1.69,    1.69,    1.69,
  1.57,    1.57,    1.57,    1.57,
  1.44,    1.44,    1.44,    1.44,
  1.37,    1.37,    1.37,    1.37,
  1.22,    1.22,    1.22,    1.22,
  1.17,    1.17,    1.17,    1.17,
  1.55,    1.55,    1.55,    1.55,
  1.99,    1.99,    1.99,    1.99,
  1.73,    1.73,    1.73,    1.73,
  1.3,     1.3,     1.3,     1.3,
  1.46,    1.46,    1.46,    1.46,
  1.14,    1.14,    1.14,    1.14,
  1.5,     1.5,     1.5,     1.5,
  1.52,    1.52,    1.52,    1.52,
  2.11,    2.11,    2.11,    2.11,
  2.47,    2.47,    2.47,    2.47,
  2.09,    2.09,    2.09,    2.09,
  2.03,    2.03,    2.03,    2.03,
  2.45,    2.45,    2.45,    2.45,
  2.7,     2.7,     2.7,     2.7,
  2.39,    2.39,    2.39,    2.39,
  2.2,     2.2,     2.2,     2.2,
  2.53,    2.53,    2.53,    2.53,
  2.37,    2.37,    2.37,    2.37,
  2.62,    2.62,    2.62,    2.62,
  2.59,    2.59,    2.59,    2.59,
  2.85,    2.85,    2.85,    2.85,
  3.09,    3.09,    3.09,    3.09,
  2.65,    2.65,    2.65,    2.65,
  2.16,    2.16,    2.16,    2.16,
  2.69,    2.69,    2.69,    2.69,
  3.49,    3.49,    3.49,    3.49,
  3.63,    3.63,    3.63,    3.63,
  3.56,    3.56,    3.56,    3.56,
  3.15,    3.15,    3.15,    3.15,
  3.76,    3.76,    3.76,    3.76,
  3.37,    3.37,    3.37,    3.37,
  3.62,    3.62,    3.62,    3.62,
  3.79,    3.79,    3.79,    3.79,
  3.57,    3.57,    3.57,    3.57,
  3.69,    3.69,    3.69,    3.69,
  3.3,     3.3,     3.3,     3.3,
  3.11,    3.11,    3.11,    3.11,
  2.75,    2.75,    2.75,    2.75,
  3.17,    3.17,    3.17,    3.17,
  2.84,    2.84,    2.84,    2.84,
  2.56,    2.56,    2.56,    2.56,
  2.49,    2.49,    2.49,    2.49,
  2.08,    2.08,    2.08,    2.08,
  2.29,    2.29,    2.29,    2.29,
  2.63,    2.63,    2.63,    2.63,
  2.67,    2.67,    2.67,    2.67,
  2.42,    2.42,    2.42,    2.42,
  2.27,    2.27,    2.27,    2.27,
  2.56,    2.56,    2.56,    2.56,
  2.29,    2.29,    2.29,    2.29,
  2.52,    2.52,    2.52,    2.52,
  2.28,    2.28,    2.28,    2.28,
  2.24,    2.24,    2.24,    2.24,
  2.17,    2.17,    2.17,    2.17,
  2.19,    2.19,    2.19,    2.19,
  2.09,    2.09,    2.09,    2.09,
  2.1,     2.1,     2.1,     2.1,
  2.07,    2.07,    2.07,    2.07,
  1.98,    1.98,    1.98,    1.98,
  1.98,    1.98,    1.98,    1.98,
  2.2,     2.2,     2.2,     2.2,
  2.41,    2.41,    2.41,    2.41,
  2.28,    2.28,    2.28,    2.28,
  2.72,    2.72,    2.72,    2.72,
  2.54,    2.54,    2.54,    2.54,
  2.68,    2.68,    2.68,    2.68,
  2.64,    2.64,    2.64,    2.64,
  2.59,    2.59,    2.59,    2.59,
  2.63,    2.63,    2.63,    2.63,
  2.21,    2.21,    2.21,    2.21,
  2.22,    2.22,    2.22,    2.22,
  1.77,    1.77,    1.77,    1.77,
  2.25,    2.25,    2.25,    2.25,
  1.71,    1.71,    1.71,    1.71,
  2.19,    2.19,    2.19,    2.19,
  2.11,    2.11,    2.11,    2.11,
  2.66,    2.66,    2.66,    2.66,
  2.76,    2.76,    2.76,    2.76,
  2.23,    2.23,    2.23,    2.23,
  2.67,    2.67,    2.67,    2.67,
  2.73,    2.73,    2.73,    2.73,
  3.3,     3.3,     3.3,     3.3,
  2.94,    2.94,    2.94,    2.94,
  2.7,     2.7,     2.7,     2.7,
  2.65,    2.65,    2.65,    2.65,
  2.43,    2.43,    2.43,    2.43,
  2.55,    2.55,    2.55,    2.55,
  2.59,    2.59,    2.59,    2.59,
  2.29,    2.29,    2.29,    2.29,
  2.48,    2.48,    2.48,    2.48,
  2.38,    2.38,    2.38,    2.38,
  2.08,    2.08,    2.08,    2.08,
  1.78,    1.78,    1.78,    1.78,
  2.1,     2.1,     2.1,     2.1,
  2.82,    2.82,    2.82,    2.82,
  3.02,    3.02,    3.02,    3.02,
  3.35,    3.35,    3.35,    3.35,
  3.26,    3.26,    3.26,    3.26,
  3.11,    3.11,    3.11,    3.11,
  2.53,    2.53,    2.53,    2.53,
  2.35,    2.35,    2.35,    2.35,
  2.43,    2.43,    2.43,    2.43,
  2.75,    2.75,    2.75,    2.75,
  2.8,     2.8,     2.8,     2.8,
  3.1,     3.1,     3.1,     3.1,
  2.97,    2.97,    2.97,    2.97,
  2.94,    2.94,    2.94,    2.94,
  2.94,    2.94,    2.94,    2.94,
  2.81,    2.81,    2.81,    2.81,
  2.89,    2.89,    2.89,    2.89,
  2.3,     2.3,     2.3,     2.3,
  2.12,    2.12,    2.12,    2.12,
  1.83,    1.83,    1.83,    1.83,
  1.82,    1.82,    1.82,    1.82,
  1.53,    1.53,    1.53,    1.53,
  1.51,    1.51,    1.51,    1.51,
  1.56,    1.56,    1.56,    1.56,
  1.08,    1.08,    1.08,    1.08,
  2.43,    2.43,    2.43,    2.43,
  2.5,     2.5,     2.5,     2.5,
  2.88,    2.88,    2.88,    2.88,
  3.16,    3.16,    3.16,    3.16,
  3.02,    3.02,    3.02,    3.02,
  3.16,    3.16,    3.16,    3.16,
  3.29,    3.29,    3.29,    3.29,
  3.08,    3.08,    3.08,    3.08,
  2.53,    2.53,    2.53,    2.53,
  2.9,     2.9,     2.9,     2.9,
  3.19,    3.19,    3.19,    3.19,
  3.57,    3.57,    3.57,    3.57,
  3.64,    3.64,    3.64,    3.64,
  3.2,     3.2,     3.2,     3.2,
  2.9,     2.9,     2.9,     2.9,
  2,       2,       2,       2,
  2.64,    2.64,    2.64,    2.64,
  2.18,    2.18,    2.18,    2.18,
  2.44,    2.44,    2.44,    2.44,
  2.32,    2.32,    2.32,    2.32,
  2.2,     2.2,     2.2,     2.2,
  2.55,    2.55,    2.55,    2.55,
  2.54,    2.54,    2.54,    2.54,
  2.53,    2.53,    2.53,    2.53,
  2.45,    2.45,    2.45,    2.45,
  2.73,    2.73,    2.73,    2.73,
  2.9,     2.9,     2.9,     2.9,
  2.52,    2.52,    2.52,    2.52,
  2.81,    2.81,    2.81,    2.81,
  2.59,    2.59,    2.59,    2.59,
  2.49,    2.49,    2.49,    2.49,
  2.44,    2.44,    2.44,    2.44,
  2.55,    2.55,    2.55,    2.55,
  2.886,   2.886,   2.886,   2.886,
  3.01,    3.01,    3.01,    3.01,
  3.113,   3.113,   3.113,   3.113,
  3.131,   3.131,   3.131,   3.131,
  3.157,   3.157,   3.157,   3.157,
  3.017,   3.017,   3.017,   3.017,
  3.208,   3.208,   3.208,   3.208,
  2.908,   2.908,   2.908,   2.908,
  2.945,   2.945,   2.945,   2.945,
  2.813,   2.813,   2.813,   2.813,
  2.69,    2.69,    2.69,    2.69,
  2.784,   2.784,   2.784,   2.784,
  2.809,   2.809,   2.809,   2.809,
  2.871,   2.871,   2.871,   2.871,
  2.76,    2.76,    2.76,    2.76,
  2.977,   2.977,   2.977,   2.977,
  2.793,   2.793,   2.793,   2.793,
  2.953,   2.953,   2.953,   2.953,
  3.215,   3.215,   3.215,   3.215,
  3.279,   3.279,   3.279,   3.279,
  3.373,   3.373,   3.373,   3.373,
  3.614,   3.614,   3.614,   3.614,
  3.583,   3.583,   3.583,   3.583,
  3.383,   3.383,   3.383,   3.383,
  3.4,     3.4,     3.4,     3.4,
  3.57,    3.57,    3.57,    3.57,
  3.477,   3.477,   3.477,   3.477,
  3.662,   3.662,   3.662,   3.662,
  3.701,   3.701,   3.701,   3.701,
  3.466,   3.466,   3.466,   3.466,
  3.47,    3.47,    3.47,    3.47,
  3.237,   3.237,   3.237,   3.237,
  2.898,   2.898,   2.898,   2.898,
  2.779,   2.779,   2.779,   2.779,
  2.61,    2.61,    2.61,    2.61,
  2.43,    2.43,    2.43,    2.43,
  2.355,   2.355,   2.355,   2.355,
  2.421,   2.421,   2.421,   2.421,
  2.621,   2.621,   2.621,   2.621,
  2.546,   2.546,   2.546,   2.546,
  2.593,   2.593,   2.593,   2.593,
  2.878,   2.878,   2.878,   2.878,
  2.945,   2.945,   2.945,   2.945,
  2.933,   2.933,   2.933,   2.933,
  2.775,   2.775,   2.775,   2.775,
  2.76,    2.76,    2.76,    2.76,
  2.706,   2.706,   2.706,   2.706,
  2.939,   2.939,   2.939,   2.939,
  2.886,   2.886,   2.886,   2.886,
  3.01,    3.01,    3.01,    3.01,
  3.113,   3.113,   3.113,   3.113,
  3.131,   3.131,   3.131,   3.131,
  3.157,   3.157,   3.157,   3.157,
  3.017,   3.017,   3.017,   3.017,
  3.208,   3.208,   3.208,   3.208,
  2.908,   2.908,   2.908,   2.908,
  2.945,   2.945,   2.945,   2.945,
  2.813,   2.813,   2.813,   2.813,
  2.69,    2.69,    2.69,    2.69,
  2.784,   2.784,   2.784,   2.784,
  2.809,   2.809,   2.809,   2.809,
  2.871,   2.871,   2.871,   2.871,
  2.76,    2.76,    2.76,    2.76,
  2.977,   2.977,   2.977,   2.977,
  2.793,   2.793,   2.793,   2.793,
  2.953,   2.953,   2.953,   2.953,
  3.215,   3.215,   3.215,   3.215,
  3.279,   3.279,   3.279,   3.279,
  3.373,   3.373,   3.373,   3.373,
  3.614,   3.614,   3.614,   3.614,
  3.583,   3.583,   3.583,   3.583,
  3.383,   3.383,   3.383,   3.383,
  3.4,     3.4,     3.4,     3.4,
  3.57,    3.57,    3.57,    3.57,
  3.477,   3.477,   3.477,   3.477,
  3.662,   3.662,   3.662,   3.662,
  3.701,   3.701,   3.701,   3.701,
  3.466,   3.466,   3.466,   3.466,
  3.47,    3.47,    3.47,    3.47,
  3.237,   3.237,   3.237,   3.237,
  2.898,   2.898,   2.898,   2.898,
  2.779,   2.779,   2.779,   2.779,
  2.61,    2.61,    2.61,    2.61,
  2.43,    2.43,    2.43,    2.43,
  2.355,   2.355,   2.355,   2.355,
  2.421,   2.421,   2.421,   2.421,
  2.621,   2.621,   2.621,   2.621,
  2.546,   2.546,   2.546,   2.546,
  2.593,   2.593,   2.593,   2.593,
  2.878,   2.878,   2.878,   2.878,
  2.945,   2.945,   2.945,   2.945,
  2.933,   2.933,   2.933,   2.933,
  2.775,   2.775,   2.775,   2.775,
  2.76,    2.76,    2.76,    2.76,
  2.706,   2.706,   2.706,   2.706,
  2.939,   2.939,   2.939,   2.939,
  2.886,   2.886,   2.886,   2.886,
  3.01,    3.01,    3.01,    3.01,
  3.113,   3.113,   3.113,   3.113,
  3.131,   3.131,   3.131,   3.131,
  3.157,   3.157,   3.157,   3.157,
  3.017,   3.017,   3.017,   3.017,
  3.208,   3.208,   3.208,   3.208,
  2.908,   2.908,   2.908,   2.908,
  2.945,   2.945,   2.945,   2.945,
  2.813,   2.813,   2.813,   2.813,
  2.69,    2.69,    2.69,    2.69,
  2.784,   2.784,   2.784,   2.784,
  2.809,   2.809,   2.809,   2.809,
  2.871,   2.871,   2.871,   2.871,
  2.76,    2.76,    2.76,    2.76,
  2.977,   2.977,   2.977,   2.977,
  2.793,   2.793,   2.793,   2.793,
  2.953,   2.953,   2.953,   2.953,
  3.215,   3.215,   3.215,   3.215,
  3.279,   3.279,   3.279,   3.279,
  3.373,   3.373,   3.373,   3.373,
  3.614,   3.614,   3.614,   3.614,
  3.583,   3.583,   3.583,   3.583,
  3.383,   3.383,   3.383,   3.383,
  3.4,     3.4,     3.4,     3.4,
  3.57,    3.57,    3.57,    3.57,
  3.477,   3.477,   3.477,   3.477,
  3.662,   3.662,   3.662,   3.662,
  3.701,   3.701,   3.701,   3.701,
  3.466,   3.466,   3.466,   3.466,
  3.47,    3.47,    3.47,    3.47,
  3.237,   3.237,   3.237,   3.237,
  2.898,   2.898,   2.898,   2.898,
  2.779,   2.779,   2.779,   2.779,
  2.61,    2.61,    2.61,    2.61,
  2.43,    2.43,    2.43,    2.43,
  2.355,   2.355,   2.355,   2.355,
  2.421,   2.421,   2.421,   2.421,
  2.621,   2.621,   2.621,   2.621,
  2.546,   2.546,   2.546,   2.546,
  2.593,   2.593,   2.593,   2.593,
  2.878,   2.878,   2.878,   2.878,
  2.945,   2.945,   2.945,   2.945,
  2.933,   2.933,   2.933,   2.933,
  2.775,   2.775,   2.775,   2.775,
  2.76,    2.76,    2.76,    2.76,
  2.706,   2.706,   2.706,   2.706,
  2.939,   2.939,   2.939,   2.939,
  2.886,   2.886,   2.886,   2.886,
  3.01,    3.01,    3.01,    3.01,
  3.113,   3.113,   3.113,   3.113,
  3.131,   3.131,   3.131,   3.131,
  3.157,   3.157,   3.157,   3.157,
  3.017,   3.017,   3.017,   3.017,
  3.208,   3.208,   3.208,   3.208,
  2.908,   2.908,   2.908,   2.908,
  2.945,   2.945,   2.945,   2.945,
  2.813,   2.813,   2.813,   2.813,
  2.69,    2.69,    2.69,    2.69,
  2.784,   2.784,   2.784,   2.784,
  2.809,   2.809,   2.809,   2.809,
  2.871,   2.871,   2.871,   2.871,
  2.76,    2.76,    2.76,    2.76,
  2.977,   2.977,   2.977,   2.977,
  2.793,   2.793,   2.793,   2.793,
  2.953,   2.953,   2.953,   2.953,
  3.215,   3.215,   3.215,   3.215,
  3.279,   3.279,   3.279,   3.279,
  3.373,   3.373,   3.373,   3.373,
  3.614,   3.614,   3.614,   3.614,
  3.583,   3.583,   3.583,   3.583,
  3.383,   3.383,   3.383,   3.383,
  3.4,     3.4,     3.4,     3.4,
  3.57,    3.57,    3.57,    3.57,
  3.477,   3.477,   3.477,   3.477,
  3.662,   3.662,   3.662,   3.662,
  3.701,   3.701,   3.701,   3.701,
  1.35,    1.35,    1.35,    1.35,
  1.29,    1.29,    1.29,    1.29,
  1.76,    1.76,    1.76,    1.76,
  2.28,    2.28,    2.28,    2.28,
  1.39,    1.39,    1.39,    1.39,
  1.79,    1.79,    1.79,    1.79,
  1.87,    1.87,    1.87,    1.87,
  2.58,    2.58,    2.58,    2.58,
  2.32,    2.32,    2.32,    2.32,
  2.3,     2.3,     2.3,     2.3,
  1.86,    1.86,    1.86,    1.86,
  1.71,    1.71,    1.71,    1.71,
  2.21,    2.21,    2.21,    2.21,
  2.19,    2.19,    2.19,    2.19,
  2.15,    2.15,    2.15,    2.15,
  1.13,    1.13,    1.13,    1.13,
  0.89,    0.89,    0.89,    0.89,
  1.18,    1.18,    1.18,    1.18,
  1.29,    1.29,    1.29,    1.29,
  0.69,    0.69,    0.69,    0.69,
  1.09,    1.09,    1.09,    1.09,
  1.47,    1.47,    1.47,    1.47,
  1.36,    1.36,    1.36,    1.36,
  1.88,    1.88,    1.88,    1.88,
  1.5,     1.5,     1.5,     1.5,
  1.25,    1.25,    1.25,    1.25,
  1.39,    1.39,    1.39,    1.39,
  1.2,     1.2,     1.2,     1.2,
  0.84,    0.84,    0.84,    0.84,
  0.58,    0.58,    0.58,    0.58,
  1.1,     1.1,     1.1,     1.1,
  1.11,    1.11,    1.11,    1.11,
  1.19,    1.19,    1.19,    1.19,
  0.81,    0.81,    0.81,    0.81,
  1.23,    1.23,    1.23,    1.23,
  1.22,    1.22,    1.22,    1.22,
  1.17,    1.17,    1.17,    1.17,
  0.9,     0.9,     0.9,     0.9,
  1.32,    1.32,    1.32,    1.32,
  1.48,    1.48,    1.48,    1.48,
  1.55,    1.55,    1.55,    1.55,
  1.42,    1.42,    1.42,    1.42,
  1.16,    1.16,    1.16,    1.16,
  0.28,    0.28,    0.28,    0.28,
  0.83,    0.83,    0.83,    0.83,
  1,       1,       1,       1,
  1.7,     1.7,     1.7,     1.7,
  1.17,    1.17,    1.17,    1.17,
  2.18,    2.18,    2.18,    2.18,
  3.21,    3.21,    3.21,    3.21,
  3.3,     3.3,     3.3,     3.3,
  2.96,    2.96,    2.96,    2.96,
  2.91,    2.91,    2.91,    2.91,
  2.48,    2.48,    2.48,    2.48,
  2.47,    2.47,    2.47,    2.47,
  0.94,    0.94,    0.94,    0.94,
  1.27,    1.27,    1.27,    1.27,
  1.94,    1.94,    1.94,    1.94,
  2.08,    2.08,    2.08,    2.08,
  2.29,    2.29,    2.29,    2.29,
  2.62,    2.62,    2.62,    2.62,
  3,       3,       3,       3,
  2.42,    2.42,    2.42,    2.42,
  2.8,     2.8,     2.8,     2.8,
  3.47,    3.47,    3.47,    3.47,
  2.96,    2.96,    2.96,    2.96,
  2.73,    2.73,    2.73,    2.73,
  3.01,    3.01,    3.01,    3.01,
  3.31,    3.31,    3.31,    3.31,
  2.28,    2.28,    2.28,    2.28,
  2.99,    2.99,    2.99,    2.99,
  2.45,    2.45,    2.45,    2.45,
  2.34,    2.34,    2.34,    2.34,
  2.3,     2.3,     2.3,     2.3,
  2.37,    2.37,    2.37,    2.37,
  2.36,    2.36,    2.36,    2.36,
  2.19,    2.19,    2.19,    2.19,
  2.72,    2.72,    2.72,    2.72,
  1.77,    1.77,    1.77,    1.77,
  1.92,    1.92,    1.92,    1.92,
  2.53,    2.53,    2.53,    2.53,
  2.28,    2.28,    2.28,    2.28,
  2.06,    2.06,    2.06,    2.06,
  2.21,    2.21,    2.21,    2.21,
  2.57,    2.57,    2.57,    2.57,
  1.72,    1.72,    1.72,    1.72,
  2.06,    2.06,    2.06,    2.06,
  2.25,    2.25,    2.25,    2.25,
  1.62,    1.62,    1.62,    1.62,
  2.09,    2.09,    2.09,    2.09,
  2.12,    2.12,    2.12,    2.12,
  2.33,    2.33,    2.33,    2.33,
  2.2,     2.2,     2.2,     2.2,
  2.13,    2.13,    2.13,    2.13,
  1.56,    1.56,    1.56,    1.56,
  1.97,    1.97,    1.97,    1.97,
  1.64,    1.64,    1.64,    1.64,
  2.24,    2.24,    2.24,    2.24,
  2.87,    2.87,    2.87,    2.87,
  2.38,    2.38,    2.38,    2.38,
  2.16,    2.16,    2.16,    2.16,
  1.86,    1.86,    1.86,    1.86,
  2.05,    2.05,    2.05,    2.05,
  2.36,    2.36,    2.36,    2.36,
  2.27,    2.27,    2.27,    2.27,
  2.18,    2.18,    2.18,    2.18,
  2.29,    2.29,    2.29,    2.29,
  2.54,    2.54,    2.54,    2.54,
  2.99,    2.99,    2.99,    2.99,
  3.35,    3.35,    3.35,    3.35,
  3.04,    3.04,    3.04,    3.04,
  2.93,    2.93,    2.93,    2.93,
  2.42,    2.42,    2.42,    2.42,
  2.25,    2.25,    2.25,    2.25,
  2.18,    2.18,    2.18,    2.18,
  2.17,    2.17,    2.17,    2.17,
  2.06,    2.06,    2.06,    2.06,
  2.15,    2.15,    2.15,    2.15,
  2.43,    2.43,    2.43,    2.43,
  2.33,    2.33,    2.33,    2.33,
  2.38,    2.38,    2.38,    2.38,
  2.4,     2.4,     2.4,     2.4,
  2.72,    2.72,    2.72,    2.72,
  2.46,    2.46,    2.46,    2.46,
  2.59,    2.59,    2.59,    2.59,
  2.26,    2.26,    2.26,    2.26,
  2.08,    2.08,    2.08,    2.08,
  2.25,    2.25,    2.25,    2.25,
  2.22,    2.22,    2.22,    2.22,
  2.53,    2.53,    2.53,    2.53,
  2.25,    2.25,    2.25,    2.25,
  2.76,    2.76,    2.76,    2.76,
  2.48,    2.48,    2.48,    2.48,
  3.21,    3.21,    3.21,    3.21,
  2.58,    2.58,    2.58,    2.58,
  2.75,    2.75,    2.75,    2.75,
  3.48,    3.48,    3.48,    3.48,
  3.2,     3.2,     3.2,     3.2,
  3,       3,       3,       3,
  3.42,    3.42,    3.42,    3.42,
  3.87,    3.87,    3.87,    3.87,
  4.13,    4.13,    4.13,    4.13,
  3.89,    3.89,    3.89,    3.89,
  3.86,    3.86,    3.86,    3.86,
  3.59,    3.59,    3.59,    3.59,
  3.94,    3.94,    3.94,    3.94,
  3.72,    3.72,    3.72,    3.72,
  3.72,    3.72,    3.72,    3.72,
  4.25,    4.25,    4.25,    4.25,
  3.59,    3.59,    3.59,    3.59,
  3.61,    3.61,    3.61,    3.61,
  3.85,    3.85,    3.85,    3.85,
  3.24,    3.24,    3.24,    3.24,
  3.93,    3.93,    3.93,    3.93,
  3.61,    3.61,    3.61,    3.61,
  4.57,    4.57,    4.57,    4.57,
  4.07,    4.07,    4.07,    4.07,
  3.39,    3.39,    3.39,    3.39,
  3.78,    3.78,    3.78,    3.78,
  3.81,    3.81,    3.81,    3.81,
  3.76,    3.76,    3.76,    3.76,
  4.09,    4.09,    4.09,    4.09,
  3.95,    3.95,    3.95,    3.95,
  4.28,    4.28,    4.28,    4.28,
  3.67,    3.67,    3.67,    3.67,
  4.05,    4.05,    4.05,    4.05,
  3.67,    3.67,    3.67,    3.67,
  3.39,    3.39,    3.39,    3.39,
  3.31,    3.31,    3.31,    3.31,
  2.47,    2.47,    2.47,    2.47,
  2.81,    2.81,    2.81,    2.81,
  2.93,    2.93,    2.93,    2.93,
  3.33,    3.33,    3.33,    3.33,
  3.49,    3.49,    3.49,    3.49,
  2.81,    2.81,    2.81,    2.81,
  2.8,     2.8,     2.8,     2.8,
  2.57,    2.57,    2.57,    2.57,
  2.84,    2.84,    2.84,    2.84,
  2.92,    2.92,    2.92,    2.92,
  3.14,    3.14,    3.14,    3.14,
  2.95,    2.95,    2.95,    2.95,
  3.43,    3.43,    3.43,    3.43,
  3.58,    3.58,    3.58,    3.58,
  3.5,     3.5,     3.5,     3.5,
  3.02,    3.02,    3.02,    3.02,
  2.42,    2.42,    2.42,    2.42,
  2.21,    2.21,    2.21,    2.21,
  2.56,    2.56,    2.56,    2.56,
  2.45,    2.45,    2.45,    2.45,
  2.39,    2.39,    2.39,    2.39,
  2.56,    2.56,    2.56,    2.56,
  2.32,    2.32,    2.32,    2.32,
  2.48,    2.48,    2.48,    2.48,
  2.77,    2.77,    2.77,    2.77,
  2.91,    2.91,    2.91,    2.91,
  2.73,    2.73,    2.73,    2.73,
  2.03,    2.03,    2.03,    2.03,
  1.98,    1.98,    1.98,    1.98,
  2.14,    2.14,    2.14,    2.14,
  2.19,    2.19,    2.19,    2.19,
  2.3,     2.3,     2.3,     2.3,
  2.83,    2.83,    2.83,    2.83,
  1.7,     1.7,     1.7,     1.7,
  1.96,    1.96,    1.96,    1.96,
  2.12,    2.12,    2.12,    2.12,
  1.98,    1.98,    1.98,    1.98,
  2.04,    2.04,    2.04,    2.04,
  2.05,    2.05,    2.05,    2.05,
  2.45,    2.45,    2.45,    2.45,
  2.38,    2.38,    2.38,    2.38,
  1.9,     1.9,     1.9,     1.9,
  1.63,    1.63,    1.63,    1.63,
  2.56,    2.56,    2.56,    2.56,
  2.42,    2.42,    2.42,    2.42,
  2.34,    2.34,    2.34,    2.34,
  2.39,    2.39,    2.39,    2.39,
  2.26,    2.26,    2.26,    2.26,
  2.41,    2.41,    2.41,    2.41,
  2.43,    2.43,    2.43,    2.43,
  2.45,    2.45,    2.45,    2.45,
  2.42,    2.42,    2.42,    2.42,
  2.4,     2.4,     2.4,     2.4,
  2.57,    2.57,    2.57,    2.57,
  2.7,     2.7,     2.7,     2.7,
  2.8,     2.8,     2.8,     2.8,
  2.52,    2.52,    2.52,    2.52,
  2.54,    2.54,    2.54,    2.54,
  2.66,    2.66,    2.66,    2.66,
  3.56,    3.56,    3.56,    3.56,
  2.98,    2.98,    2.98,    2.98,
  2.76,    2.76,    2.76,    2.76,
  3.33,    3.33,    3.33,    3.33,
  3.03,    3.03,    3.03,    3.03,
  2.94,    2.94,    2.94,    2.94,
  3.49,    3.49,    3.49,    3.49,
  3.27,    3.27,    3.27,    3.27,
  3.17,    3.17,    3.17,    3.17,
  2.75,    2.75,    2.75,    2.75,
  2.75,    2.75,    2.75,    2.75,
  2.236,   2.236,   2.236,   2.236,
  2.231,   2.231,   2.231,   2.231,
  2.354,   2.354,   2.354,   2.354,
  2.409,   2.409,   2.409,   2.409,
  2.031,   2.031,   2.031,   2.031,
  2.242,   2.242,   2.242,   2.242,
  1.957,   1.957,   1.957,   1.957,
  1.839,   1.839,   1.839,   1.839,
  2.082,   2.082,   2.082,   2.082,
  2.116,   2.116,   2.116,   2.116,
  2.25,    2.25,    2.25,    2.25,
  2.011,   2.011,   2.011,   2.011,
  2.054,   2.054,   2.054,   2.054,
  2.155,   2.155,   2.155,   2.155,
  1.973,   1.973,   1.973,   1.973,
  2.144,   2.144,   2.144,   2.144,
  2.228,   2.228,   2.228,   2.228,
  2.162,   2.162,   2.162,   2.162,
  2.147,   2.147,   2.147,   2.147,
  2.129,   2.129,   2.129,   2.129,
  2.105,   2.105,   2.105,   2.105,
  2.11,    2.11,    2.11,    2.11,
  2.034,   2.034,   2.034,   2.034,
  2.004,   2.004,   2.004,   2.004,
  1.897,   1.897,   1.897,   1.897,
  1.997,   1.997,   1.997,   1.997,
  1.989,   1.989,   1.989,   1.989,
  2.026,   2.026,   2.026,   2.026,
  1.957,   1.957,   1.957,   1.957,
  2.049,   2.049,   2.049,   2.049,
  2.22,    2.22,    2.22,    2.22,
  1.998,   1.998,   1.998,   1.998,
  2.088,   2.088,   2.088,   2.088,
  2.044,   2.044,   2.044,   2.044,
  2.15,    2.15,    2.15,    2.15,
  2.173,   2.173,   2.173,   2.173,
  2.019,   2.019,   2.019,   2.019,
  2.365,   2.365,   2.365,   2.365,
  2.468,   2.468,   2.468,   2.468,
  2.415,   2.415,   2.415,   2.415,
  2.497,   2.497,   2.497,   2.497,
  2.353,   2.353,   2.353,   2.353,
  2.37,    2.37,    2.37,    2.37,
  2.327,   2.327,   2.327,   2.327,
  2.538,   2.538,   2.538,   2.538,
  2.627,   2.627,   2.627,   2.627,
  2.41,    2.41,    2.41,    2.41,
  2.197,   2.197,   2.197,   2.197,
  2.236,   2.236,   2.236,   2.236,
  2.231,   2.231,   2.231,   2.231,
  2.354,   2.354,   2.354,   2.354,
  2.409,   2.409,   2.409,   2.409,
  2.031,   2.031,   2.031,   2.031,
  2.242,   2.242,   2.242,   2.242,
  1.957,   1.957,   1.957,   1.957,
  1.839,   1.839,   1.839,   1.839,
  2.082,   2.082,   2.082,   2.082,
  2.116,   2.116,   2.116,   2.116,
  2.25,    2.25,    2.25,    2.25,
  2.011,   2.011,   2.011,   2.011,
  2.054,   2.054,   2.054,   2.054,
  2.155,   2.155,   2.155,   2.155,
  1.973,   1.973,   1.973,   1.973,
  2.144,   2.144,   2.144,   2.144,
  2.228,   2.228,   2.228,   2.228,
  2.162,   2.162,   2.162,   2.162,
  2.147,   2.147,   2.147,   2.147,
  2.129,   2.129,   2.129,   2.129,
  2.105,   2.105,   2.105,   2.105,
  2.11,    2.11,    2.11,    2.11,
  2.034,   2.034,   2.034,   2.034,
  2.004,   2.004,   2.004,   2.004,
  1.897,   1.897,   1.897,   1.897,
  1.997,   1.997,   1.997,   1.997,
  1.989,   1.989,   1.989,   1.989,
  2.026,   2.026,   2.026,   2.026,
  1.957,   1.957,   1.957,   1.957,
  2.049,   2.049,   2.049,   2.049,
  2.22,    2.22,    2.22,    2.22,
  1.998,   1.998,   1.998,   1.998,
  2.088,   2.088,   2.088,   2.088,
  2.044,   2.044,   2.044,   2.044,
  2.15,    2.15,    2.15,    2.15,
  2.173,   2.173,   2.173,   2.173,
  2.019,   2.019,   2.019,   2.019,
  2.365,   2.365,   2.365,   2.365,
  2.468,   2.468,   2.468,   2.468,
  2.415,   2.415,   2.415,   2.415,
  2.497,   2.497,   2.497,   2.497,
  2.353,   2.353,   2.353,   2.353,
  2.37,    2.37,    2.37,    2.37,
  2.327,   2.327,   2.327,   2.327,
  2.538,   2.538,   2.538,   2.538,
  2.627,   2.627,   2.627,   2.627,
  2.41,    2.41,    2.41,    2.41,
  2.197,   2.197,   2.197,   2.197,
  2.236,   2.236,   2.236,   2.236,
  2.231,   2.231,   2.231,   2.231,
  2.354,   2.354,   2.354,   2.354,
  2.409,   2.409,   2.409,   2.409,
  2.031,   2.031,   2.031,   2.031,
  2.242,   2.242,   2.242,   2.242,
  1.957,   1.957,   1.957,   1.957,
  1.839,   1.839,   1.839,   1.839,
  2.082,   2.082,   2.082,   2.082,
  2.116,   2.116,   2.116,   2.116,
  2.25,    2.25,    2.25,    2.25,
  2.011,   2.011,   2.011,   2.011,
  2.054,   2.054,   2.054,   2.054,
  2.155,   2.155,   2.155,   2.155,
  1.973,   1.973,   1.973,   1.973,
  2.144,   2.144,   2.144,   2.144,
  2.228,   2.228,   2.228,   2.228,
  2.162,   2.162,   2.162,   2.162,
  2.147,   2.147,   2.147,   2.147,
  2.129,   2.129,   2.129,   2.129,
  2.105,   2.105,   2.105,   2.105,
  2.11,    2.11,    2.11,    2.11,
  2.034,   2.034,   2.034,   2.034,
  2.004,   2.004,   2.004,   2.004,
  1.897,   1.897,   1.897,   1.897,
  1.997,   1.997,   1.997,   1.997,
  1.989,   1.989,   1.989,   1.989,
  2.026,   2.026,   2.026,   2.026,
  1.957,   1.957,   1.957,   1.957,
  2.049,   2.049,   2.049,   2.049,
  2.22,    2.22,    2.22,    2.22,
  1.998,   1.998,   1.998,   1.998,
  2.088,   2.088,   2.088,   2.088,
  2.044,   2.044,   2.044,   2.044,
  2.15,    2.15,    2.15,    2.15,
  2.173,   2.173,   2.173,   2.173,
  2.019,   2.019,   2.019,   2.019,
  2.365,   2.365,   2.365,   2.365,
  2.468,   2.468,   2.468,   2.468,
  2.415,   2.415,   2.415,   2.415,
  2.497,   2.497,   2.497,   2.497,
  2.353,   2.353,   2.353,   2.353,
  2.37,    2.37,    2.37,    2.37,
  2.327,   2.327,   2.327,   2.327,
  2.538,   2.538,   2.538,   2.538,
  2.627,   2.627,   2.627,   2.627,
  2.41,    2.41,    2.41,    2.41,
  2.197,   2.197,   2.197,   2.197,
  2.236,   2.236,   2.236,   2.236,
  2.231,   2.231,   2.231,   2.231,
  2.354,   2.354,   2.354,   2.354,
  2.409,   2.409,   2.409,   2.409,
  2.031,   2.031,   2.031,   2.031,
  2.242,   2.242,   2.242,   2.242,
  1.957,   1.957,   1.957,   1.957,
  1.839,   1.839,   1.839,   1.839,
  2.082,   2.082,   2.082,   2.082,
  2.116,   2.116,   2.116,   2.116,
  2.25,    2.25,    2.25,    2.25,
  2.011,   2.011,   2.011,   2.011,
  2.054,   2.054,   2.054,   2.054,
  2.155,   2.155,   2.155,   2.155,
  1.973,   1.973,   1.973,   1.973,
  2.144,   2.144,   2.144,   2.144,
  2.228,   2.228,   2.228,   2.228,
  2.162,   2.162,   2.162,   2.162,
  2.147,   2.147,   2.147,   2.147,
  2.129,   2.129,   2.129,   2.129,
  2.105,   2.105,   2.105,   2.105,
  2.11,    2.11,    2.11,    2.11,
  2.034,   2.034,   2.034,   2.034,
  2.004,   2.004,   2.004,   2.004,
  1.897,   1.897,   1.897,   1.897,
  1.997,   1.997,   1.997,   1.997,
  1.989,   1.989,   1.989,   1.989,
  2.026,   2.026,   2.026,   2.026,
  1.957,   1.957,   1.957,   1.957,
  2.049,   2.049,   2.049,   2.049,
  2.22,    2.22,    2.22,    2.22,
  1.998,   1.998,   1.998,   1.998,
  2.088,   2.088,   2.088,   2.088,
  2.044,   2.044,   2.044,   2.044,
  2.15,    2.15,    2.15,    2.15,
  2.173,   2.173,   2.173,   2.173,
  2.019,   2.019,   2.019,   2.019,
  2.365,   2.365,   2.365,   2.365,
  2.468,   2.468,   2.468,   2.468,
  2.415,   2.415,   2.415,   2.415,
  2.497,   2.497,   2.497,   2.497,
  2.353,   2.353,   2.353,   2.353,
  2.37,    2.37,    2.37,    2.37,
  2.327,   2.327,   2.327,   2.327,
  2.538,   2.538,   2.538,   2.538,
  2.627,   2.627,   2.627,   2.627,
  2.41,    2.41,    2.41,    2.41,
  2.197,   2.197,   2.197,   2.197,
  2.236,   2.236,   2.236,   2.236,
  2.231,   2.231,   2.231,   2.231,
  2.354,   2.354,   2.354,   2.354,
  2.409,   2.409,   2.409,   2.409,
  2.031,   2.031,   2.031,   2.031,
  4.62,    4.62,    4.62,    4.62,
  4.3,     4.3,     4.3,     4.3,
  3.09,    3.09,    3.09,    3.09,
  3.45,    3.45,    3.45,    3.45,
  3.61,    3.61,    3.61,    3.61,
  3.96,    3.96,    3.96,    3.96,
  3.17,    3.17,    3.17,    3.17,
  2.66,    2.66,    2.66,    2.66,
  3.56,    3.56,    3.56,    3.56,
  2.99,    2.99,    2.99,    2.99,
  3,       3,       3,       3,
  3.05,    3.05,    3.05,    3.05,
  2.8,     2.8,     2.8,     2.8,
  2.51,    2.51,    2.51,    2.51,
  2.63,    2.63,    2.63,    2.63,
  2.12,    2.12,    2.12,    2.12,
  1.77,    1.77,    1.77,    1.77,
  2.18,    2.18,    2.18,    2.18,
  1.33,    1.33,    1.33,    1.33,
  1.55,    1.55,    1.55,    1.55,
  1.65,    1.65,    1.65,    1.65,
  1.23,    1.23,    1.23,    1.23,
  1.49,    1.49,    1.49,    1.49,
  1.03,    1.03,    1.03,    1.03,
  1.27,    1.27,    1.27,    1.27,
  1.02,    1.02,    1.02,    1.02,
  1.22,    1.22,    1.22,    1.22,
  1.39,    1.39,    1.39,    1.39,
  0.41,    0.41,    0.41,    0.41,
  0.48,    0.48,    0.48,    0.48,
  0.88,    0.88,    0.88,    0.88,
  0.89,    0.89,    0.89,    0.89,
  1.8,     1.8,     1.8,     1.8,
  1.78,    1.78,    1.78,    1.78,
  1.89,    1.89,    1.89,    1.89,
  2.45,    2.45,    2.45,    2.45,
  2.27,    2.27,    2.27,    2.27,
  2.82,    2.82,    2.82,    2.82,
  2.19,    2.19,    2.19,    2.19,
  2.83,    2.83,    2.83,    2.83,
  2.86,    2.86,    2.86,    2.86,
  2.49,    2.49,    2.49,    2.49,
  1.61,    1.61,    1.61,    1.61,
  1.97,    1.97,    1.97,    1.97,
  1.93,    1.93,    1.93,    1.93,
  2.29,    2.29,    2.29,    2.29,
  2.55,    2.55,    2.55,    2.55,
  1.95,    1.95,    1.95,    1.95,
  2.11,    2.11,    2.11,    2.11,
  0.44,    0.44,    0.44,    0.44,
  1.57,    1.57,    1.57,    1.57,
  1.89,    1.89,    1.89,    1.89,
  2.27,    2.27,    2.27,    2.27,
  2.42,    2.42,    2.42,    2.42,
  2.51,    2.51,    2.51,    2.51,
  2.24,    2.24,    2.24,    2.24,
  1.9,     1.9,     1.9,     1.9,
  1.41,    1.41,    1.41,    1.41,
  2.32,    2.32,    2.32,    2.32,
  2.41,    2.41,    2.41,    2.41,
  2.08,    2.08,    2.08,    2.08,
  1.99,    1.99,    1.99,    1.99,
  2.3,     2.3,     2.3,     2.3,
  2.3,     2.3,     2.3,     2.3,
  2.5,     2.5,     2.5,     2.5,
  2.47,    2.47,    2.47,    2.47,
  3.04,    3.04,    3.04,    3.04,
  2.56,    2.56,    2.56,    2.56,
  3.21,    3.21,    3.21,    3.21,
  3.51,    3.51,    3.51,    3.51,
  3.59,    3.59,    3.59,    3.59,
  3.7,     3.7,     3.7,     3.7,
  3.66,    3.66,    3.66,    3.66,
  4.28,    4.28,    4.28,    4.28,
  3.59,    3.59,    3.59,    3.59,
  3.45,    3.45,    3.45,    3.45,
  3.15,    3.15,    3.15,    3.15,
  3.63,    3.63,    3.63,    3.63,
  3.57,    3.57,    3.57,    3.57,
  3.01,    3.01,    3.01,    3.01,
  3.78,    3.78,    3.78,    3.78,
  4.38,    4.38,    4.38,    4.38,
  4.75,    4.75,    4.75,    4.75,
  4.08,    4.08,    4.08,    4.08,
  3.81,    3.81,    3.81,    3.81,
  3.87,    3.87,    3.87,    3.87,
  4.02,    4.02,    4.02,    4.02,
  3.89,    3.89,    3.89,    3.89,
  4.31,    4.31,    4.31,    4.31,
  4.3,     4.3,     4.3,     4.3,
  3.74,    3.74,    3.74,    3.74,
  3.73,    3.73,    3.73,    3.73,
  4.15,    4.15,    4.15,    4.15,
  3.95,    3.95,    3.95,    3.95,
  3.96,    3.96,    3.96,    3.96,
  3.32,    3.32,    3.32,    3.32,
  3.86,    3.86,    3.86,    3.86,
  3.28,    3.28,    3.28,    3.28,
  3.35,    3.35,    3.35,    3.35,
  3.33,    3.33,    3.33,    3.33,
  3.13,    3.13,    3.13,    3.13,
  2.38,    2.38,    2.38,    2.38,
  2.15,    2.15,    2.15,    2.15,
  1.83,    1.83,    1.83,    1.83,
  1.83,    1.83,    1.83,    1.83,
  1.58,    1.58,    1.58,    1.58,
  1.39,    1.39,    1.39,    1.39,
  1.39,    1.39,    1.39,    1.39,
  1.51,    1.51,    1.51,    1.51,
  1.4,     1.4,     1.4,     1.4,
  1.1,     1.1,     1.1,     1.1,
  1.16,    1.16,    1.16,    1.16,
  0.37,    0.37,    0.37,    0.37,
  1.38,    1.38,    1.38,    1.38,
  1.67,    1.67,    1.67,    1.67,
  1.34,    1.34,    1.34,    1.34,
  1.04,    1.04,    1.04,    1.04,
  0.94,    0.94,    0.94,    0.94,
  0.59,    0.59,    0.59,    0.59,
  0.71,    0.71,    0.71,    0.71,
  0.18,    0.18,    0.18,    0.18,
  0.4,     0.4,     0.4,     0.4,
  0.82,    0.82,    0.82,    0.82,
  1.38,    1.38,    1.38,    1.38,
  1.78,    1.78,    1.78,    1.78,
  1.14,    1.14,    1.14,    1.14,
  1.59,    1.59,    1.59,    1.59,
  0.69,    0.69,    0.69,    0.69,
  0.99,    0.99,    0.99,    0.99,
  1.16,    1.16,    1.16,    1.16,
  1.04,    1.04,    1.04,    1.04,
  1.58,    1.58,    1.58,    1.58,
  1.28,    1.28,    1.28,    1.28,
  1.43,    1.43,    1.43,    1.43,
  1.68,    1.68,    1.68,    1.68,
  2.01,    2.01,    2.01,    2.01,
  1.7,     1.7,     1.7,     1.7,
  1.99,    1.99,    1.99,    1.99,
  1.78,    1.78,    1.78,    1.78,
  1.84,    1.84,    1.84,    1.84,
  1.91,    1.91,    1.91,    1.91,
  1.86,    1.86,    1.86,    1.86,
  1.64,    1.64,    1.64,    1.64,
  1.2,     1.2,     1.2,     1.2,
  1.22,    1.22,    1.22,    1.22,
  1.55,    1.55,    1.55,    1.55,
  1.43,    1.43,    1.43,    1.43,
  1.42,    1.42,    1.42,    1.42,
  1.6,     1.6,     1.6,     1.6,
  2.06,    2.06,    2.06,    2.06,
  1.99,    1.99,    1.99,    1.99,
  1.7,     1.7,     1.7,     1.7,
  1.69,    1.69,    1.69,    1.69,
  1.68,    1.68,    1.68,    1.68,
  2,       2,       2,       2,
  2.18,    2.18,    2.18,    2.18,
  2.6,     2.6,     2.6,     2.6,
  3.07,    3.07,    3.07,    3.07,
  2.78,    2.78,    2.78,    2.78,
  2.36,    2.36,    2.36,    2.36,
  2.1,     2.1,     2.1,     2.1,
  1.3,     1.3,     1.3,     1.3,
  1.7,     1.7,     1.7,     1.7,
  2.1,     2.1,     2.1,     2.1,
  2.46,    2.46,    2.46,    2.46,
  2.38,    2.38,    2.38,    2.38,
  2.72,    2.72,    2.72,    2.72,
  2.47,    2.47,    2.47,    2.47,
  2.86,    2.86,    2.86,    2.86,
  3.06,    3.06,    3.06,    3.06,
  3.04,    3.04,    3.04,    3.04,
  3.27,    3.27,    3.27,    3.27,
  3.02,    3.02,    3.02,    3.02,
  3.86,    3.86,    3.86,    3.86,
  3.69,    3.69,    3.69,    3.69,
  3.62,    3.62,    3.62,    3.62,
  3.96,    3.96,    3.96,    3.96,
  4.09,    4.09,    4.09,    4.09,
  3.55,    3.55,    3.55,    3.55,
  3.2,     3.2,     3.2,     3.2,
  3.68,    3.68,    3.68,    3.68,
  3.05,    3.05,    3.05,    3.05,
  2.9,     2.9,     2.9,     2.9,
  2.65,    2.65,    2.65,    2.65,
  2.81,    2.81,    2.81,    2.81,
  2.85,    2.85,    2.85,    2.85,
  1.84,    1.84,    1.84,    1.84,
  2.3,     2.3,     2.3,     2.3,
  1.92,    1.92,    1.92,    1.92,
  1.66,    1.66,    1.66,    1.66,
  1.59,    1.59,    1.59,    1.59,
  0.84,    0.84,    0.84,    0.84,
  0.79,    0.79,    0.79,    0.79,
  0.92,    0.92,    0.92,    0.92,
  0.12,    0.12,    0.12,    0.12,
  0.48,    0.48,    0.48,    0.48,
  0.64,    0.64,    0.64,    0.64,
  0.29,    0.29,    0.29,    0.29,
  0.22,    0.22,    0.22,    0.22,
  0.18,    0.18,    0.18,    0.18,
  0.46,    0.46,    0.46,    0.46,
  0.34,    0.34,    0.34,    0.34,
  0.9,     0.9,     0.9,     0.9,
  1.11,    1.11,    1.11,    1.11,
  0.81,    0.81,    0.81,    0.81,
  0.59,    0.59,    0.59,    0.59,
  0.58,    0.58,    0.58,    0.58,
  1.11,    1.11,    1.11,    1.11,
  1.87,    1.87,    1.87,    1.87,
  1.39,    1.39,    1.39,    1.39,
  0.7,     0.7,     0.7,     0.7,
  0.48,    0.48,    0.48,    0.48,
  0.55,    0.55,    0.55,    0.55,
  1.15,    1.15,    1.15,    1.15,
  0.92,    0.92,    0.92,    0.92,
  1.09,    1.09,    1.09,    1.09,
  1.39,    1.39,    1.39,    1.39,
  1.58,    1.58,    1.58,    1.58,
  1.11,    1.11,    1.11,    1.11,
  0.92,    0.92,    0.92,    0.92,
  1.06,    1.06,    1.06,    1.06,
  1.42,    1.42,    1.42,    1.42,
  1.64,    1.64,    1.64,    1.64,
  0.91,    0.91,    0.91,    0.91,
  0.88,    0.88,    0.88,    0.88,
  0.98,    0.98,    0.98,    0.98,
  1.25,    1.25,    1.25,    1.25,
  0.92,    0.92,    0.92,    0.92,
  0.98,    0.98,    0.98,    0.98,
  1.4,     1.4,     1.4,     1.4,
  1.24,    1.24,    1.24,    1.24,
  1.29,    1.29,    1.29,    1.29,
  1.44,    1.44,    1.44,    1.44,
  0.97,    0.97,    0.97,    0.97,
  1.49,    1.49,    1.49,    1.49,
  1.17,    1.17,    1.17,    1.17,
  1.32,    1.32,    1.32,    1.32,
  1.25,    1.25,    1.25,    1.25,
  1.04,    1.04,    1.04,    1.04,
  0.64,    0.64,    0.64,    0.64,
  0.3,     0.3,     0.3,     0.3,
  0.94,    0.94,    0.94,    0.94,
  0.4,     0.4,     0.4,     0.4,
  0.69,    0.69,    0.69,    0.69,
  0.81,    0.81,    0.81,    0.81,
  0.58,    0.58,    0.58,    0.58,
  0.55,    0.55,    0.55,    0.55,
  1.1,     1.1,     1.1,     1.1,
  1.06,    1.06,    1.06,    1.06,
  1.24,    1.24,    1.24,    1.24,
  1.08,    1.08,    1.08,    1.08,
  1.26,    1.26,    1.26,    1.26,
  1.27,    1.27,    1.27,    1.27,
  1.33,    1.33,    1.33,    1.33,
  1.14,    1.14,    1.14,    1.14,
  0.91,    0.91,    0.91,    0.91,
  0.89,    0.89,    0.89,    0.89,
  0.72,    0.72,    0.72,    0.72,
  0.17,    0.17,    0.17,    0.17,
  0.38,    0.38,    0.38,    0.38,
  0.77,    0.77,    0.77,    0.77,
  1.1,     1.1,     1.1,     1.1,
  0.62,    0.62,    0.62,    0.62,
  0.37,    0.37,    0.37,    0.37,
  0.6,     0.6,     0.6,     0.6,
  0.99,    0.99,    0.99,    0.99,
  0.97,    0.97,    0.97,    0.97,
  0.8,     0.8,     0.8,     0.8,
  0.9,     0.9,     0.9,     0.9,
  0.8,     0.8,     0.8,     0.8,
  0.59,    0.59,    0.59,    0.59,
  0.3,     0.3,     0.3,     0.3,
  0.68,    0.68,    0.68,    0.68,
  0.95,    0.95,    0.95,    0.95,
  0.69,    0.69,    0.69,    0.69,
  0.91,    0.91,    0.91,    0.91,
  0.36,    0.36,    0.36,    0.36,
  0.48,    0.48,    0.48,    0.48,
  0.42,    0.42,    0.42,    0.42,
  1.13,    1.13,    1.13,    1.13,
  1.46,    1.46,    1.46,    1.46,
  0.1,     0.1,     0.1,     0.1,
  0.75,    0.75,    0.75,    0.75,
  0.96,    0.96,    0.96,    0.96,
  1.14,    1.14,    1.14,    1.14,
  1.23,    1.23,    1.23,    1.23,
  1.4,     1.4,     1.4,     1.4,
  1.5,     1.5,     1.5,     1.5,
  1.08,    1.08,    1.08,    1.08,
  0.71,    0.71,    0.71,    0.71,
  0.63,    0.63,    0.63,    0.63,
  1.16,    1.16,    1.16,    1.16,
  1.29,    1.29,    1.29,    1.29,
  1.87,    1.87,    1.87,    1.87,
  1.92,    1.92,    1.92,    1.92,
  1.76,    1.76,    1.76,    1.76,
  1.87,    1.87,    1.87,    1.87,
  1.77,    1.77,    1.77,    1.77,
  1.89,    1.89,    1.89,    1.89,
  2.09,    2.09,    2.09,    2.09,
  1.92,    1.92,    1.92,    1.92,
  1.86,    1.86,    1.86,    1.86,
  1.86,    1.86,    1.86,    1.86,
  1.99,    1.99,    1.99,    1.99,
  1.79,    1.79,    1.79,    1.79,
  1.46,    1.46,    1.46,    1.46,
  1.86,    1.86,    1.86,    1.86,
  1.96,    1.96,    1.96,    1.96,
  1.76,    1.76,    1.76,    1.76,
  1.66,    1.66,    1.66,    1.66,
  1.69,    1.69,    1.69,    1.69,
  2.09,    2.09,    2.09,    2.09,
  2.15,    2.15,    2.15,    2.15,
  2.39,    2.39,    2.39,    2.39,
  2.35,    2.35,    2.35,    2.35,
  2.23,    2.23,    2.23,    2.23,
  2.29,    2.29,    2.29,    2.29,
  2.67,    2.67,    2.67,    2.67,
  2.97,    2.97,    2.97,    2.97,
  2.97,    2.97,    2.97,    2.97,
  3.2,     3.2,     3.2,     3.2,
  3.6,     3.6,     3.6,     3.6,
  3.58,    3.58,    3.58,    3.58,
  3.79,    3.79,    3.79,    3.79,
  4.39,    4.39,    4.39,    4.39,
  4.04,    4.04,    4.04,    4.04,
  3.86,    3.86,    3.86,    3.86,
  4.59,    4.59,    4.59,    4.59,
  4.52,    4.52,    4.52,    4.52,
  4.45,    4.45,    4.45,    4.45,
  5.12,    5.12,    5.12,    5.12,
  4.89,    4.89,    4.89,    4.89,
  5.5,     5.5,     5.5,     5.5,
  5.36,    5.36,    5.36,    5.36,
  5.23,    5.23,    5.23,    5.23,
  5.14,    5.14,    5.14,    5.14,
  4.97,    4.97,    4.97,    4.97,
  4.99,    4.99,    4.99,    4.99,
  5.43,    5.43,    5.43,    5.43,
  6.11,    6.11,    6.11,    6.11,
  5.74,    5.74,    5.74,    5.74,
  5.56,    5.56,    5.56,    5.56,
  4.36,    4.36,    4.36,    4.36,
  4.75,    4.75,    4.75,    4.75,
  4.52,    4.52,    4.52,    4.52,
  5.04,    5.04,    5.04,    5.04,
  5.2,     5.2,     5.2,     5.2,
  4.74,    4.74,    4.74,    4.74,
  4.13,    4.13,    4.13,    4.13,
  3.91,    3.91,    3.91,    3.91,
  4.06,    4.06,    4.06,    4.06,
  4.29,    4.29,    4.29,    4.29,
  4.33,    4.33,    4.33,    4.33,
  4.01,    4.01,    4.01,    4.01,
  3.3,     3.3,     3.3,     3.3,
  3.03,    3.03,    3.03,    3.03,
  2.68,    2.68,    2.68,    2.68,
  3.25,    3.25,    3.25,    3.25,
  3.51,    3.51,    3.51,    3.51,
  3.12,    3.12,    3.12,    3.12,
  3.36,    3.36,    3.36,    3.36,
  3.22,    3.22,    3.22,    3.22,
  2.87,    2.87,    2.87,    2.87,
  2.43,    2.43,    2.43,    2.43,
  2.82,    2.82,    2.82,    2.82,
  2.65,    2.65,    2.65,    2.65,
  2.19,    2.19,    2.19,    2.19,
  2.85,    2.85,    2.85,    2.85,
  3.24,    3.24,    3.24,    3.24,
  4.62,    4.62,    4.62,    4.62,
  4.75,    4.75,    4.75,    4.75,
  4.38,    4.38,    4.38,    4.38,
  4.66,    4.66,    4.66,    4.66,
  4.93,    4.93,    4.93,    4.93,
  4.83,    4.83,    4.83,    4.83,
  5.84,    5.84,    5.84,    5.84,
  5.35,    5.35,    5.35,    5.35,
  5.86,    5.86,    5.86,    5.86,
  5.45,    5.45,    5.45,    5.45,
  5,       5,       5,       5,
  5.73,    5.73,    5.73,    5.73,
  4.8,     4.8,     4.8,     4.8,
  4.88,    4.88,    4.88,    4.88,
  4.81,    4.81,    4.81,    4.81,
  3.64,    3.64,    3.64,    3.64,
  3.86,    3.86,    3.86,    3.86,
  2.87,    2.87,    2.87,    2.87,
  3,       3,       3,       3,
  4.14,    4.14,    4.14,    4.14,
  4.79,    4.79,    4.79,    4.79,
  6.25,    6.25,    6.25,    6.25,
  5.72,    5.72,    5.72,    5.72,
  6.39,    6.39,    6.39,    6.39,
  6.82,    6.82,    6.82,    6.82,
  6.71,    6.71,    6.71,    6.71,
  6.52,    6.52,    6.52,    6.52,
  7.26,    7.26,    7.26,    7.26,
  7.73,    7.73,    7.73,    7.73,
  7.47,    7.47,    7.47,    7.47,
  7.16,    7.16,    7.16,    7.16,
  7.44,    7.44,    7.44,    7.44,
  6.2,     6.2,     6.2,     6.2,
  9.92,    9.92,    9.92,    9.92,
  9.35,    9.35,    9.35,    9.35,
  8.47,    8.47,    8.47,    8.47,
  7.92,    7.92,    7.92,    7.92,
  7.06,    7.06,    7.06,    7.06,
  4.67,    4.67,    4.67,    4.67,
  5.06,    5.06,    5.06,    5.06,
  4.6,     4.6,     4.6,     4.6,
  5.27,    5.27,    5.27,    5.27,
  5.49,    5.49,    5.49,    5.49,
  5.84,    5.84,    5.84,    5.84,
  6.15,    6.15,    6.15,    6.15,
  5.45,    5.45,    5.45,    5.45,
  5.74,    5.74,    5.74,    5.74,
  5.22,    5.22,    5.22,    5.22,
  6.32,    6.32,    6.32,    6.32,
  6.63,    6.63,    6.63,    6.63,
  6.97,    6.97,    6.97,    6.97,
  6.78,    6.78,    6.78,    6.78,
  6.92,    6.92,    6.92,    6.92,
  7.35,    7.35,    7.35,    7.35,
  7.14,    7.14,    7.14,    7.14,
  6.79,    6.79,    6.79,    6.79,
  6.45,    6.45,    6.45,    6.45,
  6.75,    6.75,    6.75,    6.75,
  7.11,    7.11,    7.11,    7.11,
  6.87,    6.87,    6.87,    6.87,
  6.41,    6.41,    6.41,    6.41,
  6.12,    6.12,    6.12,    6.12,
  6.26,    6.26,    6.26,    6.26,
  6.29,    6.29,    6.29,    6.29,
  5.96,    5.96,    5.96,    5.96,
  6.38,    6.38,    6.38,    6.38,
  5.25,    5.25,    5.25,    5.25,
  5.09,    5.09,    5.09,    5.09,
  5.62,    5.62,    5.62,    5.62,
  4.97,    4.97,    4.97,    4.97,
  4.46,    4.46,    4.46,    4.46,
  4.78,    4.78,    4.78,    4.78,
  4.55,    4.55,    4.55,    4.55,
  4,       4,       4,       4,
  3.83,    3.83,    3.83,    3.83,
  3.74,    3.74,    3.74,    3.74,
  3.35,    3.35,    3.35,    3.35,
  3.26,    3.26,    3.26,    3.26,
  3.06,    3.06,    3.06,    3.06,
  3.82,    3.82,    3.82,    3.82,
  3.8,     3.8,     3.8,     3.8,
  3.5,     3.5,     3.5,     3.5,
  3.35,    3.35,    3.35,    3.35,
  3.15,    3.15,    3.15,    3.15,
  3.18,    3.18,    3.18,    3.18,
  3.26,    3.26,    3.26,    3.26,
  3.97,    3.97,    3.97,    3.97,
  4.25,    4.25,    4.25,    4.25,
  3.88,    3.88,    3.88,    3.88,
  4.4,     4.4,     4.4,     4.4,
  4.12,    4.12,    4.12,    4.12,
  3.86,    3.86,    3.86,    3.86,
  3.66,    3.66,    3.66,    3.66,
  3.8,     3.8,     3.8,     3.8,
  4.36,    4.36,    4.36,    4.36,
  4.78,    4.78,    4.78,    4.78,
  5.26,    5.26,    5.26,    5.26,
  4.9,     4.9,     4.9,     4.9,
  5.84,    5.84,    5.84,    5.84,
  5.36,    5.36,    5.36,    5.36,
  4.72,    4.72,    4.72,    4.72,
  5.25,    5.25,    5.25,    5.25,
  5.44,    5.44,    5.44,    5.44,
  5.05,    5.05,    5.05,    5.05,
  5.34,    5.34,    5.34,    5.34,
  5.21,    5.21,    5.21,    5.21,
  4.68,    4.68,    4.68,    4.68,
  5.1,     5.1,     5.1,     5.1,
  4.23,    4.23,    4.23,    4.23,
  3.81,    3.81,    3.81,    3.81,
  4.73,    4.73,    4.73,    4.73,
  4.07,    4.07,    4.07,    4.07,
  3.92,    3.92,    3.92,    3.92,
  3.37,    3.37,    3.37,    3.37,
  3.48,    3.48,    3.48,    3.48,
  3.76,    3.76,    3.76,    3.76,
  2.63,    2.63,    2.63,    2.63,
  2.39,    2.39,    2.39,    2.39,
  2.64,    2.64,    2.64,    2.64,
  2.93,    2.93,    2.93,    2.93,
  2.27,    2.27,    2.27,    2.27,
  2.65,    2.65,    2.65,    2.65,
  2.6,     2.6,     2.6,     2.6,
  2.98,    2.98,    2.98,    2.98,
  2.97,    2.97,    2.97,    2.97,
  2.84,    2.84,    2.84,    2.84,
  2.66,    2.66,    2.66,    2.66,
  2.85,    2.85,    2.85,    2.85,
  2.77,    2.77,    2.77,    2.77,
  2.3,     2.3,     2.3,     2.3,
  2.11,    2.11,    2.11,    2.11,
  1.76,    1.76,    1.76,    1.76,
  1.76,    1.76,    1.76,    1.76,
  1.69,    1.69,    1.69,    1.69,
  1.9,     1.9,     1.9,     1.9,
  1.87,    1.87,    1.87,    1.87,
  1.38,    1.38,    1.38,    1.38,
  1.82,    1.82,    1.82,    1.82,
  1.69,    1.69,    1.69,    1.69,
  1.48,    1.48,    1.48,    1.48,
  1.49,    1.49,    1.49,    1.49,
  1.43,    1.43,    1.43,    1.43,
  2.05,    2.05,    2.05,    2.05,
  2.54,    2.54,    2.54,    2.54,
  3.04,    3.04,    3.04,    3.04,
  3.47,    3.47,    3.47,    3.47,
  3.33,    3.33,    3.33,    3.33,
  3.14,    3.14,    3.14,    3.14,
  2.75,    2.75,    2.75,    2.75,
  2.82,    2.82,    2.82,    2.82,
  3.37,    3.37,    3.37,    3.37,
  3.27,    3.27,    3.27,    3.27,
  2.67,    2.67,    2.67,    2.67,
  2.75,    2.75,    2.75,    2.75,
  4.23,    4.23,    4.23,    4.23,
  4.09,    4.09,    4.09,    4.09,
  4.04,    4.04,    4.04,    4.04,
  4.05,    4.05,    4.05,    4.05,
  4.03,    4.03,    4.03,    4.03,
  3.55,    3.55,    3.55,    3.55,
  3.01,    3.01,    3.01,    3.01,
  2.89,    2.89,    2.89,    2.89,
  2.45,    2.45,    2.45,    2.45,
  2.36,    2.36,    2.36,    2.36,
  2.36,    2.36,    2.36,    2.36,
  2.28,    2.28,    2.28,    2.28,
  1.95,    1.95,    1.95,    1.95,
  1.87,    1.87,    1.87,    1.87,
  2,       2,       2,       2,
  2.06,    2.06,    2.06,    2.06,
  1.95,    1.95,    1.95,    1.95,
  1.82,    1.82,    1.82,    1.82,
  1.88,    1.88,    1.88,    1.88,
  1.69,    1.69,    1.69,    1.69,
  0.99,    0.99,    0.99,    0.99,
  1.53,    1.53,    1.53,    1.53,
  2.01,    2.01,    2.01,    2.01,
  2.19,    2.19,    2.19,    2.19,
  2.13,    2.13,    2.13,    2.13,
  1.79,    1.79,    1.79,    1.79,
  1.97,    1.97,    1.97,    1.97,
  2.16,    2.16,    2.16,    2.16,
  2.08,    2.08,    2.08,    2.08,
  2.03,    2.03,    2.03,    2.03,
  1.59,    1.59,    1.59,    1.59,
  1.62,    1.62,    1.62,    1.62,
  2.15,    2.15,    2.15,    2.15,
  1.92,    1.92,    1.92,    1.92,
  1.82,    1.82,    1.82,    1.82,
  1.62,    1.62,    1.62,    1.62,
  1.63,    1.63,    1.63,    1.63,
  2.9,     2.9,     2.9,     2.9,
  3.24,    3.24,    3.24,    3.24,
  3.8,     3.8,     3.8,     3.8,
  3.55,    3.55,    3.55,    3.55,
  3.11,    3.11,    3.11,    3.11,
  3.2,     3.2,     3.2,     3.2,
  3.02,    3.02,    3.02,    3.02,
  2.92,    2.92,    2.92,    2.92,
  3.29,    3.29,    3.29,    3.29,
  2.82,    2.82,    2.82,    2.82,
  2.58,    2.58,    2.58,    2.58,
  3.1,     3.1,     3.1,     3.1,
  3.01,    3.01,    3.01,    3.01,
  2.58,    2.58,    2.58,    2.58,
  2.43,    2.43,    2.43,    2.43,
  2.72,    2.72,    2.72,    2.72,
  2.6,     2.6,     2.6,     2.6,
  2.32,    2.32,    2.32,    2.32,
  2.12,    2.12,    2.12,    2.12,
  1.64,    1.64,    1.64,    1.64,
  1.97,    1.97,    1.97,    1.97,
  1.96,    1.96,    1.96,    1.96,
  2.28,    2.28,    2.28,    2.28,
  1.65,    1.65,    1.65,    1.65,
  1.27,    1.27,    1.27,    1.27,
  1.68,    1.68,    1.68,    1.68,
  2.33,    2.33,    2.33,    2.33,
  2.63,    2.63,    2.63,    2.63,
  2.62,    2.62,    2.62,    2.62,
  2.81,    2.81,    2.81,    2.81,
  2.53,    2.53,    2.53,    2.53,
  2.7,     2.7,     2.7,     2.7,
  2.82,    2.82,    2.82,    2.82,
  2.58,    2.58,    2.58,    2.58,
  2.37,    2.37,    2.37,    2.37,
  2.54,    2.54,    2.54,    2.54,
  2.37,    2.37,    2.37,    2.37,
  2.1,     2.1,     2.1,     2.1,
  1.72,    1.72,    1.72,    1.72,
  2.33,    2.33,    2.33,    2.33,
  2.42,    2.42,    2.42,    2.42,
  2.33,    2.33,    2.33,    2.33,
  2.28,    2.28,    2.28,    2.28,
  2.21,    2.21,    2.21,    2.21,
  2.28,    2.28,    2.28,    2.28,
  1.84,    1.84,    1.84,    1.84,
  1.36,    1.36,    1.36,    1.36,
  1.22,    1.22,    1.22,    1.22,
  1.79,    1.79,    1.79,    1.79,
  2.3,     2.3,     2.3,     2.3,
  2.55,    2.55,    2.55,    2.55,
  2.59,    2.59,    2.59,    2.59,
  2.7,     2.7,     2.7,     2.7,
  2.97,    2.97,    2.97,    2.97,
  3.39,    3.39,    3.39,    3.39,
  2.82,    2.82,    2.82,    2.82,
  2.45,    2.45,    2.45,    2.45,
  3.04,    3.04,    3.04,    3.04,
  2.6,     2.6,     2.6,     2.6,
  3.36,    3.36,    3.36,    3.36,
  3.42,    3.42,    3.42,    3.42,
  2.47,    2.47,    2.47,    2.47,
  2.74,    2.74,    2.74,    2.74,
  3.01,    3.01,    3.01,    3.01,
  3,       3,       3,       3,
  2.95,    2.95,    2.95,    2.95,
  2.93,    2.93,    2.93,    2.93,
  2.2,     2.2,     2.2,     2.2,
  2.1,     2.1,     2.1,     2.1,
  2.15,    2.15,    2.15,    2.15,
  2.39,    2.39,    2.39,    2.39,
  2.34,    2.34,    2.34,    2.34,
  2.22,    2.22,    2.22,    2.22,
  2.21,    2.21,    2.21,    2.21,
  2.2,     2.2,     2.2,     2.2,
  1.71,    1.71,    1.71,    1.71,
  0.82,    0.82,    0.82,    0.82,
  0.58,    0.58,    0.58,    0.58,
  0.62,    0.62,    0.62,    0.62,
  0.36,    0.36,    0.36,    0.36,
  0.68,    0.68,    0.68,    0.68,
  0.42,    0.42,    0.42,    0.42,
  0.92,    0.92,    0.92,    0.92,
  0.68,    0.68,    0.68,    0.68,
  1.09,    1.09,    1.09,    1.09,
  1.07,    1.07,    1.07,    1.07,
  1.69,    1.69,    1.69,    1.69,
  2.16,    2.16,    2.16,    2.16,
  2.35,    2.35,    2.35,    2.35,
  2.23,    2.23,    2.23,    2.23,
  2.06,    2.06,    2.06,    2.06,
  1.95,    1.95,    1.95,    1.95,
  1.75,    1.75,    1.75,    1.75,
  1.41,    1.41,    1.41,    1.41,
  0.65,    0.65,    0.65,    0.65,
  0.45,    0.45,    0.45,    0.45,
  0.51,    0.51,    0.51,    0.51,
  0.6,     0.6,     0.6,     0.6,
  0.84,    0.84,    0.84,    0.84,
  1.16,    1.16,    1.16,    1.16,
  1.17,    1.17,    1.17,    1.17,
  1.78,    1.78,    1.78,    1.78,
  1.85,    1.85,    1.85,    1.85,
  2.16,    2.16,    2.16,    2.16,
  1.94,    1.94,    1.94,    1.94,
  2.44,    2.44,    2.44,    2.44,
  2.46,    2.46,    2.46,    2.46,
  1.99,    1.99,    1.99,    1.99,
  1.54,    1.54,    1.54,    1.54,
  1.77,    1.77,    1.77,    1.77,
  2.31,    2.31,    2.31,    2.31,
  1.87,    1.87,    1.87,    1.87,
  0.96,    0.96,    0.96,    0.96,
  1.47,    1.47,    1.47,    1.47,
  1.99,    1.99,    1.99,    1.99,
  1.51,    1.51,    1.51,    1.51,
  1.18,    1.18,    1.18,    1.18,
  1.57,    1.57,    1.57,    1.57,
  2.01,    2.01,    2.01,    2.01,
  1.87,    1.87,    1.87,    1.87,
  1.36,    1.36,    1.36,    1.36,
  1.33,    1.33,    1.33,    1.33,
  1.39,    1.39,    1.39,    1.39,
  1.91,    1.91,    1.91,    1.91,
  1.82,    1.82,    1.82,    1.82,
  1.66,    1.66,    1.66,    1.66,
  1.93,    1.93,    1.93,    1.93,
  1.72,    1.72,    1.72,    1.72,
  1.23,    1.23,    1.23,    1.23,
  1.47,    1.47,    1.47,    1.47,
  1.67,    1.67,    1.67,    1.67,
  1.5,     1.5,     1.5,     1.5,
  1.66,    1.66,    1.66,    1.66,
  2.04,    2.04,    2.04,    2.04,
  2.04,    2.04,    2.04,    2.04,
  1.72,    1.72,    1.72,    1.72,
  1.85,    1.85,    1.85,    1.85,
  2.52,    2.52,    2.52,    2.52,
  2.27,    2.27,    2.27,    2.27,
  1.4,     1.4,     1.4,     1.4,
  1.2,     1.2,     1.2,     1.2,
  2.3,     2.3,     2.3,     2.3,
  2.25,    2.25,    2.25,    2.25,
  2.9,     2.9,     2.9,     2.9,
  3.08,    3.08,    3.08,    3.08,
  4.57,    4.57,    4.57,    4.57,
  4.79,    4.79,    4.79,    4.79,
  4.76,    4.76,    4.76,    4.76,
  4.9,     4.9,     4.9,     4.9,
  5.98,    5.98,    5.98,    5.98,
  5.46,    5.46,    5.46,    5.46,
  5.95,    5.95,    5.95,    5.95,
  6.49,    6.49,    6.49,    6.49,
  5.81,    5.81,    5.81,    5.81,
  4.39,    4.39,    4.39,    4.39,
  6.19,    6.19,    6.19,    6.19,
  6.26,    6.26,    6.26,    6.26,
  7.01,    7.01,    7.01,    7.01,
  6.79,    6.79,    6.79,    6.79,
  6.97,    6.97,    6.97,    6.97,
  6.52,    6.52,    6.52,    6.52,
  5.87,    5.87,    5.87,    5.87,
  5.66,    5.66,    5.66,    5.66,
  5.87,    5.87,    5.87,    5.87,
  4.08,    4.08,    4.08,    4.08,
  3.45,    3.45,    3.45,    3.45,
  2.83,    2.83,    2.83,    2.83,
  2.78,    2.78,    2.78,    2.78,
  2.34,    2.34,    2.34,    2.34,
  2.47,    2.47,    2.47,    2.47,
  2.43,    2.43,    2.43,    2.43,
  2.34,    2.34,    2.34,    2.34,
  2.56,    2.56,    2.56,    2.56,
  2.38,    2.38,    2.38,    2.38,
  2.943,   2.943,   2.943,   2.943,
  3.46,    3.46,    3.46,    3.46,
  4.98,    4.98,    4.98,    4.98,
  4.88,    4.88,    4.88,    4.88,
  4.58,    4.58,    4.58,    4.58,
  4.22,    4.22,    4.22,    4.22,
  3.58,    3.58,    3.58,    3.58,
  4.6,     4.6,     4.6,     4.6,
  3.5,     3.5,     3.5,     3.5,
  4.03,    4.03,    4.03,    4.03,
  3.72,    3.72,    3.72,    3.72,
  3.14,    3.14,    3.14,    3.14,
  3.44,    3.44,    3.44,    3.44,
  3.54,    3.54,    3.54,    3.54,
  4.19,    4.19,    4.19,    4.19,
  4.73,    4.73,    4.73,    4.73,
  3.61,    3.61,    3.61,    3.61,
  4.54,    4.54,    4.54,    4.54,
  5.28,    5.28,    5.28,    5.28,
  4.96,    4.96,    4.96,    4.96,
  4.3,     4.3,     4.3,     4.3,
  4.56,    4.56,    4.56,    4.56,
  4.63,    4.63,    4.63,    4.63,
  5.71,    5.71,    5.71,    5.71,
  4.63,    4.63,    4.63,    4.63,
  5.95,    5.95,    5.95,    5.95,
  5.55,    5.55,    5.55,    5.55,
  5.34,    5.34,    5.34,    5.34,
  5.67,    5.67,    5.67,    5.67,
  5.86,    5.86,    5.86,    5.86,
  4.8,     4.8,     4.8,     4.8,
  5.42,    5.42,    5.42,    5.42,
  5.28,    5.28,    5.28,    5.28,
  5.07,    5.07,    5.07,    5.07,
  4.65,    4.65,    4.65,    4.65,
  4.59,    4.59,    4.59,    4.59,
  4.83,    4.83,    4.83,    4.83,
  3.79,    3.79,    3.79,    3.79,
  3.24,    3.24,    3.24,    3.24,
  2.6,     2.6,     2.6,     2.6,
  2.55,    2.55,    2.55,    2.55,
  2.09,    2.09,    2.09,    2.09,
  1.42,    1.42,    1.42,    1.42,
  1.69,    1.69,    1.69,    1.69,
  1.96,    1.96,    1.96,    1.96,
  2.12,    2.12,    2.12,    2.12,
  1.91,    1.91,    1.91,    1.91,
  2.6,     2.6,     2.6,     2.6,
  2.48,    2.48,    2.48,    2.48,
  2.83,    2.83,    2.83,    2.83,
  3.03,    3.03,    3.03,    3.03,
  3.44,    3.44,    3.44,    3.44,
  4.2,     4.2,     4.2,     4.2,
  4.19,    4.19,    4.19,    4.19,
  4.33,    4.33,    4.33,    4.33,
  4.4,     4.4,     4.4,     4.4,
  3.79,    3.79,    3.79,    3.79,
  3.42,    3.42,    3.42,    3.42,
  3.48,    3.48,    3.48,    3.48,
  3.4,     3.4,     3.4,     3.4,
  3.5,     3.5,     3.5,     3.5,
  4.38,    4.38,    4.38,    4.38,
  4.45,    4.45,    4.45,    4.45,
  4.51,    4.51,    4.51,    4.51,
  4.84,    4.84,    4.84,    4.84,
  4.91,    4.91,    4.91,    4.91,
  5.14,    5.14,    5.14,    5.14,
  4.98,    4.98,    4.98,    4.98,
  4.94,    4.94,    4.94,    4.94,
  5.14,    5.14,    5.14,    5.14,
  5.01,    5.01,    5.01,    5.01,
  4.86,    4.86,    4.86,    4.86,
  4.99,    4.99,    4.99,    4.99,
  4.94,    4.94,    4.94,    4.94,
  5.31,    5.31,    5.31,    5.31,
  5.7,     5.7,     5.7,     5.7,
  5.66,    5.66,    5.66,    5.66,
  5.68,    5.68,    5.68,    5.68,
  5.41,    5.41,    5.41,    5.41,
  5.51,    5.51,    5.51,    5.51,
  5.99,    5.99,    5.99,    5.99,
  5.72,    5.72,    5.72,    5.72,
  5.33,    5.33,    5.33,    5.33,
  5.88,    5.88,    5.88,    5.88,
  6.15,    6.15,    6.15,    6.15,
  6.5,     6.5,     6.5,     6.5,
  5.37,    5.37,    5.37,    5.37,
  5.77,    5.77,    5.77,    5.77,
  6.19,    6.19,    6.19,    6.19,
  6.83,    6.83,    6.83,    6.83,
  6.66,    6.66,    6.66,    6.66,
  5.84,    5.84,    5.84,    5.84,
  6.89,    6.89,    6.89,    6.89,
  7.12,    7.12,    7.12,    7.12,
  5.48,    5.48,    5.48,    5.48,
  4.64,    4.64,    4.64,    4.64,
  5.4,     5.4,     5.4,     5.4,
  4.21,    4.21,    4.21,    4.21,
  4,       4,       4,       4,
  2.93,    2.93,    2.93,    2.93,
  3.122,   3.122,   3.122,   3.122,
  3.025,   3.025,   3.025,   3.025,
  3.26,    3.26,    3.26,    3.26,
  3.2,     3.2,     3.2,     3.2,
  2.85,    2.85,    2.85,    2.85,
  1.94,    1.94,    1.94,    1.94,
  1.7,     1.7,     1.7,     1.7,
  1.8,     1.8,     1.8,     1.8,
  2.07,    2.07,    2.07,    2.07,
  2.08,    2.08,    2.08,    2.08,
  1.92,    1.92,    1.92,    1.92,
  1.47,    1.47,    1.47,    1.47,
  1.85,    1.85,    1.85,    1.85,
  2.38,    2.38,    2.38,    2.38,
  2.7,     2.7,     2.7,     2.7,
  2.84,    2.84,    2.84,    2.84,
  3.26,    3.26,    3.26,    3.26,
  2.57,    2.57,    2.57,    2.57,
  2.5,     2.5,     2.5,     2.5,
  3.25,    3.25,    3.25,    3.25,
  3.39,    3.39,    3.39,    3.39,
  3.49,    3.49,    3.49,    3.49,
  3.17,    3.17,    3.17,    3.17,
  3.91,    3.91,    3.91,    3.91,
  3.49,    3.49,    3.49,    3.49,
  3.9,     3.9,     3.9,     3.9,
  4.12,    4.12,    4.12,    4.12,
  4.09,    4.09,    4.09,    4.09,
  4.3,     4.3,     4.3,     4.3,
  4.57,    4.57,    4.57,    4.57,
  3.86,    3.86,    3.86,    3.86,
  3.96,    3.96,    3.96,    3.96,
  2.91,    2.91,    2.91,    2.91,
  2.61,    2.61,    2.61,    2.61,
  2.25,    2.25,    2.25,    2.25,
  1.92,    1.92,    1.92,    1.92,
  1.61,    1.61,    1.61,    1.61,
  2.26,    2.26,    2.26,    2.26,
  2.49,    2.49,    2.49,    2.49,
  2.23,    2.23,    2.23,    2.23,
  1.89,    1.89,    1.89,    1.89,
  2.03,    2.03,    2.03,    2.03,
  2.12,    2.12,    2.12,    2.12,
  1.62,    1.62,    1.62,    1.62,
  1.58,    1.58,    1.58,    1.58,
  1.09,    1.09,    1.09,    1.09,
  1.18,    1.18,    1.18,    1.18,
  1.03,    1.03,    1.03,    1.03,
  0.73,    0.73,    0.73,    0.73,
  1.25,    1.25,    1.25,    1.25,
  1.31,    1.31,    1.31,    1.31,
  1.61,    1.61,    1.61,    1.61,
  0.96,    0.96,    0.96,    0.96,
  1.02,    1.02,    1.02,    1.02,
  1.68,    1.68,    1.68,    1.68,
  2.1,     2.1,     2.1,     2.1,
  1.64,    1.64,    1.64,    1.64,
  1.56,    1.56,    1.56,    1.56,
  1.72,    1.72,    1.72,    1.72,
  1.3,     1.3,     1.3,     1.3,
  1.09,    1.09,    1.09,    1.09,
  1.75,    1.75,    1.75,    1.75,
  1.78,    1.78,    1.78,    1.78,
  0.74,    0.74,    0.74,    0.74,
  2.06,    2.06,    2.06,    2.06,
  2.23,    2.23,    2.23,    2.23,
  2.05,    2.05,    2.05,    2.05,
  2.29,    2.29,    2.29,    2.29,
  2.3,     2.3,     2.3,     2.3,
  2.08,    2.08,    2.08,    2.08,
  1.45,    1.45,    1.45,    1.45,
  1.25,    1.25,    1.25,    1.25,
  1.87,    1.87,    1.87,    1.87,
  1.74,    1.74,    1.74,    1.74,
  1.59,    1.59,    1.59,    1.59,
  1.44,    1.44,    1.44,    1.44,
  2.16,    2.16,    2.16,    2.16,
  2.54,    2.54,    2.54,    2.54,
  2.34,    2.34,    2.34,    2.34,
  2.1,     2.1,     2.1,     2.1,
  2.31,    2.31,    2.31,    2.31,
  2.22,    2.22,    2.22,    2.22,
  1.95,    1.95,    1.95,    1.95,
  2.17,    2.17,    2.17,    2.17,
  2.28,    2.28,    2.28,    2.28,
  2.47,    2.47,    2.47,    2.47,
  2.75,    2.75,    2.75,    2.75,
  2.85,    2.85,    2.85,    2.85,
  2.94,    2.94,    2.94,    2.94,
  2.58,    2.58,    2.58,    2.58,
  2.38,    2.38,    2.38,    2.38,
  2.17,    2.17,    2.17,    2.17,
  2.54,    2.54,    2.54,    2.54,
  2.68,    2.68,    2.68,    2.68,
  2.64,    2.64,    2.64,    2.64,
  2.95,    2.95,    2.95,    2.95,
  3.04,    3.04,    3.04,    3.04,
  3.01,    3.01,    3.01,    3.01,
  2.98,    2.98,    2.98,    2.98,
  2.66,    2.66,    2.66,    2.66,
  2.35,    2.35,    2.35,    2.35,
  1.97,    1.97,    1.97,    1.97,
  2.24,    2.24,    2.24,    2.24,
  2.24,    2.24,    2.24,    2.24,
  2.22,    2.22,    2.22,    2.22,
  2.23,    2.23,    2.23,    2.23,
  2.07,    2.07,    2.07,    2.07,
  1.93,    1.93,    1.93,    1.93,
  2.16,    2.16,    2.16,    2.16,
  2.8,     2.8,     2.8,     2.8,
  2.85,    2.85,    2.85,    2.85,
  2.82,    2.82,    2.82,    2.82,
  3,       3,       3,       3,
  2.66,    2.66,    2.66,    2.66,
  1.95,    1.95,    1.95,    1.95,
  2.35,    2.35,    2.35,    2.35,
  1.75,    1.75,    1.75,    1.75,
  2.08,    2.08,    2.08,    2.08,
  2.07,    2.07,    2.07,    2.07,
  2,       2,       2,       2,
  1.55,    1.55,    1.55,    1.55,
  1.69,    1.69,    1.69,    1.69,
  1.88,    1.88,    1.88,    1.88,
  2.18,    2.18,    2.18,    2.18,
  2.72,    2.72,    2.72,    2.72,
  3.02,    3.02,    3.02,    3.02,
  2.31,    2.31,    2.31,    2.31,
  2.19,    2.19,    2.19,    2.19,
  2.87,    2.87,    2.87,    2.87,
  2.19,    2.19,    2.19,    2.19,
  1.97,    1.97,    1.97,    1.97,
  2.46,    2.46,    2.46,    2.46,
  2.43,    2.43,    2.43,    2.43,
  2.61,    2.61,    2.61,    2.61,
  2.68,    2.68,    2.68,    2.68,
  2.72,    2.72,    2.72,    2.72,
  2.76,    2.76,    2.76,    2.76,
  2.41,    2.41,    2.41,    2.41,
  2.49,    2.49,    2.49,    2.49,
  2.49,    2.49,    2.49,    2.49,
  2.51,    2.51,    2.51,    2.51,
  2.38,    2.38,    2.38,    2.38,
  2.36,    2.36,    2.36,    2.36,
  2.51,    2.51,    2.51,    2.51,
  2.42,    2.42,    2.42,    2.42,
  2.38,    2.38,    2.38,    2.38,
  2.27,    2.27,    2.27,    2.27,
  2.37,    2.37,    2.37,    2.37,
  2.13,    2.13,    2.13,    2.13,
  2.09,    2.09,    2.09,    2.09,
  2.19,    2.19,    2.19,    2.19,
  2.06,    2.06,    2.06,    2.06,
  2.12,    2.12,    2.12,    2.12,
  2.13,    2.13,    2.13,    2.13,
  2.27,    2.27,    2.27,    2.27,
  1.53,    1.53,    1.53,    1.53,
  1.58,    1.58,    1.58,    1.58,
  1.66,    1.66,    1.66,    1.66,
  1.5,     1.5,     1.5,     1.5,
  1,       1,       1,       1,
  0.88,    0.88,    0.88,    0.88,
  1.28,    1.28,    1.28,    1.28,
  0.8,     0.8,     0.8,     0.8,
  0.98,    0.98,    0.98,    0.98,
  0.79,    0.79,    0.79,    0.79,
  0.91,    0.91,    0.91,    0.91,
  1.69,    1.69,    1.69,    1.69,
  1.43,    1.43,    1.43,    1.43,
  1.67,    1.67,    1.67,    1.67,
  1.82,    1.82,    1.82,    1.82,
  1.87,    1.87,    1.87,    1.87,
  1.53,    1.53,    1.53,    1.53,
  1.23,    1.23,    1.23,    1.23,
  1.63,    1.63,    1.63,    1.63,
  2.17,    2.17,    2.17,    2.17,
  2.79,    2.79,    2.79,    2.79,
  2.28,    2.28,    2.28,    2.28,
  1.87,    1.87,    1.87,    1.87,
  2.25,    2.25,    2.25,    2.25,
  2.17,    2.17,    2.17,    2.17,
  2.24,    2.24,    2.24,    2.24,
  1.96,    1.96,    1.96,    1.96,
  2.13,    2.13,    2.13,    2.13,
  2.01,    2.01,    2.01,    2.01,
  2,       2,       2,       2,
  2.49,    2.49,    2.49,    2.49,
  1.93,    1.93,    1.93,    1.93,
  0.96,    0.96,    0.96,    0.96,
  0.76,    0.76,    0.76,    0.76,
  0.68,    0.68,    0.68,    0.68,
  2.096,   2.096,   2.096,   2.096,
  1.49,    1.49,    1.49,    1.49,
  1.2,     1.2,     1.2,     1.2,
  1.22,    1.22,    1.22,    1.22,
  1.53,    1.53,    1.53,    1.53,
  1.05,    1.05,    1.05,    1.05,
  1.38,    1.38,    1.38,    1.38,
  1.76,    1.76,    1.76,    1.76,
  1.63,    1.63,    1.63,    1.63,
  0.91,    0.91,    0.91,    0.91,
  1.27,    1.27,    1.27,    1.27,
  0.72,    0.72,    0.72,    0.72,
  0.58,    0.58,    0.58,    0.58,
  0.46,    0.46,    0.46,    0.46,
  0.5,     0.5,     0.5,     0.5,
  0.53,    0.53,    0.53,    0.53,
  1.07,    1.07,    1.07,    1.07,
  1.5,     1.5,     1.5,     1.5,
  1.58,    1.58,    1.58,    1.58,
  1.43,    1.43,    1.43,    1.43,
  1.73,    1.73,    1.73,    1.73,
  1.73,    1.73,    1.73,    1.73,
  2.19,    2.19,    2.19,    2.19,
  2.89,    2.89,    2.89,    2.89,
  2.92,    2.92,    2.92,    2.92,
  3.16,    3.16,    3.16,    3.16,
  3.28,    3.28,    3.28,    3.28,
  2.951,   2.951,   2.951,   2.951,
  2.758,   2.758,   2.758,   2.758,
  2.99,    2.99,    2.99,    2.99,
  2.87,    2.87,    2.87,    2.87,
  3.26,    3.26,    3.26,    3.26,
  3.18,    3.18,    3.18,    3.18,
  3.33,    3.33,    3.33,    3.33,
  2.6,     2.6,     2.6,     2.6,
  2.39,    2.39,    2.39,    2.39,
  2.04,    2.04,    2.04,    2.04,
  1.91,    1.91,    1.91,    1.91,
  2.16,    2.16,    2.16,    2.16,
  1.89,    1.89,    1.89,    1.89,
  1.89,    1.89,    1.89,    1.89,
  2.21,    2.21,    2.21,    2.21,
  2.08,    2.08,    2.08,    2.08,
  2,       2,       2,       2,
  2.14,    2.14,    2.14,    2.14,
  2.08,    2.08,    2.08,    2.08,
  2.23,    2.23,    2.23,    2.23,
  2.28,    2.28,    2.28,    2.28,
  2.096,   2.096,   2.096,   2.096,
  2.66,    2.66,    2.66,    2.66,
  2.46,    2.46,    2.46,    2.46,
  2.2,     2.2,     2.2,     2.2,
  1.99,    1.99,    1.99,    1.99,
  2.22,    2.22,    2.22,    2.22,
  2.2,     2.2,     2.2,     2.2,
  2.2,     2.2,     2.2,     2.2,
  2.56,    2.56,    2.56,    2.56,
  2.69,    2.69,    2.69,    2.69,
  2.78,    2.78,    2.78,    2.78,
  2.98,    2.98,    2.98,    2.98,
  2.87,    2.87,    2.87,    2.87,
  3.12,    3.12,    3.12,    3.12,
  3.6,     3.6,     3.6,     3.6,
  4.46,    4.46,    4.46,    4.46,
  5.49,    5.49,    5.49,    5.49,
  5.6,     5.6,     5.6,     5.6,
  5.84,    5.84,    5.84,    5.84,
  6.6,     6.6,     6.6,     6.6,
  2.699,   2.699,   2.699,   2.699,
  2.472,   2.472,   2.472,   2.472,
  2.788,   2.788,   2.788,   2.788,
  2.717,   2.717,   2.717,   2.717,
  2.65,    2.65,    2.65,    2.65,
  2.658,   2.658,   2.658,   2.658,
  2.913,   2.913,   2.913,   2.913,
  2.951,   2.951,   2.951,   2.951,
  2.758,   2.758,   2.758,   2.758,
  3.027,   3.027,   3.027,   3.027,
  3.261,   3.261,   3.261,   3.261,
  3.397,   3.397,   3.397,   3.397,
  3.241,   3.241,   3.241,   3.241,
  3.291,   3.291,   3.291,   3.291,
  2.969,   2.969,   2.969,   2.969,
  2.818,   2.818,   2.818,   2.818,
  2.595,   2.595,   2.595,   2.595,
  2.324,   2.324,   2.324,   2.324,
  2.327,   2.327,   2.327,   2.327,
  2.148,   2.148,   2.148,   2.148,
  2.04,    2.04,    2.04,    2.04,
  2.22,    2.22,    2.22,    2.22,
  2.112,   2.112,   2.112,   2.112,
  1.974,   1.974,   1.974,   1.974,
  2.04,    2.04,    2.04,    2.04,
  1.902,   1.902,   1.902,   1.902,
  1.937,   1.937,   1.937,   1.937,
  1.982,   1.982,   1.982,   1.982,
  2.096,   2.096,   2.096,   2.096,
  2.008,   2.008,   2.008,   2.008,
  2.02,    2.02,    2.02,    2.02,
  1.989,   1.989,   1.989,   1.989,
  1.891,   1.891,   1.891,   1.891,
  1.921,   1.921,   1.921,   1.921,
  1.884,   1.884,   1.884,   1.884,
  1.834,   1.834,   1.834,   1.834,
  1.925,   1.925,   1.925,   1.925,
  1.809,   1.809,   1.809,   1.809,
  1.685,   1.685,   1.685,   1.685,
  1.535,   1.535,   1.535,   1.535,
  1.555,   1.555,   1.555,   1.555,
  1.534,   1.534,   1.534,   1.534,
  1.805,   1.805,   1.805,   1.805,
  2.165,   2.165,   2.165,   2.165,
  2.55,    2.55,    2.55,    2.55,
  2.78,    2.78,    2.78,    2.78,
  2.763,   2.763,   2.763,   2.763,
  2.97,    2.97,    2.97,    2.97,
  2.699,   2.699,   2.699,   2.699,
  2.472,   2.472,   2.472,   2.472,
  2.788,   2.788,   2.788,   2.788,
  2.717,   2.717,   2.717,   2.717,
  2.65,    2.65,    2.65,    2.65,
  2.658,   2.658,   2.658,   2.658,
  2.913,   2.913,   2.913,   2.913,
  2.951,   2.951,   2.951,   2.951,
  2.758,   2.758,   2.758,   2.758,
  3.027,   3.027,   3.027,   3.027,
  3.261,   3.261,   3.261,   3.261,
  3.397,   3.397,   3.397,   3.397,
  3.241,   3.241,   3.241,   3.241,
  3.291,   3.291,   3.291,   3.291,
  2.969,   2.969,   2.969,   2.969,
  2.818,   2.818,   2.818,   2.818,
  2.595,   2.595,   2.595,   2.595,
  2.324,   2.324,   2.324,   2.324,
  2.327,   2.327,   2.327,   2.327,
  2.148,   2.148,   2.148,   2.148,
  2.04,    2.04,    2.04,    2.04,
  2.22,    2.22,    2.22,    2.22,
  2.112,   2.112,   2.112,   2.112,
  1.974,   1.974,   1.974,   1.974,
  2.04,    2.04,    2.04,    2.04,
  1.902,   1.902,   1.902,   1.902,
  1.937,   1.937,   1.937,   1.937,
  1.982,   1.982,   1.982,   1.982,
  2.096,   2.096,   2.096,   2.096,
  2.008,   2.008,   2.008,   2.008,
  2.02,    2.02,    2.02,    2.02,
  1.989,   1.989,   1.989,   1.989,
  1.891,   1.891,   1.891,   1.891,
  1.921,   1.921,   1.921,   1.921,
  1.884,   1.884,   1.884,   1.884,
  1.834,   1.834,   1.834,   1.834,
  1.925,   1.925,   1.925,   1.925,
  1.809,   1.809,   1.809,   1.809,
  1.685,   1.685,   1.685,   1.685,
  1.535,   1.535,   1.535,   1.535,
  1.555,   1.555,   1.555,   1.555,
  1.534,   1.534,   1.534,   1.534,
  1.805,   1.805,   1.805,   1.805,
  2.165,   2.165,   2.165,   2.165,
  2.55,    2.55,    2.55,    2.55,
  2.78,    2.78,    2.78,    2.78,
  2.763,   2.763,   2.763,   2.763,
  2.97,    2.97,    2.97,    2.97,
  2.699,   2.699,   2.699,   2.699,
  2.472,   2.472,   2.472,   2.472,
  2.788,   2.788,   2.788,   2.788,
  2.717,   2.717,   2.717,   2.717,
  2.65,    2.65,    2.65,    2.65,
  2.658,   2.658,   2.658,   2.658,
  2.913,   2.913,   2.913,   2.913,
  2.951,   2.951,   2.951,   2.951,
  2.758,   2.758,   2.758,   2.758,
  3.027,   3.027,   3.027,   3.027,
  3.261,   3.261,   3.261,   3.261,
  3.397,   3.397,   3.397,   3.397,
  3.241,   3.241,   3.241,   3.241,
  3.291,   3.291,   3.291,   3.291,
  2.969,   2.969,   2.969,   2.969,
  2.818,   2.818,   2.818,   2.818,
  2.595,   2.595,   2.595,   2.595,
  2.324,   2.324,   2.324,   2.324,
  2.327,   2.327,   2.327,   2.327,
  2.148,   2.148,   2.148,   2.148,
  2.04,    2.04,    2.04,    2.04,
  2.22,    2.22,    2.22,    2.22,
  2.112,   2.112,   2.112,   2.112,
  1.974,   1.974,   1.974,   1.974,
  2.04,    2.04,    2.04,    2.04,
  1.902,   1.902,   1.902,   1.902,
  1.937,   1.937,   1.937,   1.937,
  1.982,   1.982,   1.982,   1.982,
  2.096,   2.096,   2.096,   2.096,
  2.008,   2.008,   2.008,   2.008,
  2.02,    2.02,    2.02,    2.02,
  1.989,   1.989,   1.989,   1.989,
  1.891,   1.891,   1.891,   1.891,
  1.921,   1.921,   1.921,   1.921,
  1.884,   1.884,   1.884,   1.884,
  1.834,   1.834,   1.834,   1.834,
  1.925,   1.925,   1.925,   1.925,
  1.809,   1.809,   1.809,   1.809,
  1.685,   1.685,   1.685,   1.685,
  1.535,   1.535,   1.535,   1.535,
  1.555,   1.555,   1.555,   1.555,
  1.534,   1.534,   1.534,   1.534,
  1.805,   1.805,   1.805,   1.805,
  2.165,   2.165,   2.165,   2.165,
  2.55,    2.55,    2.55,    2.55,
  2.78,    2.78,    2.78,    2.78,
  2.763,   2.763,   2.763,   2.763,
  2.97,    2.97,    2.97,    2.97,
  2.699,   2.699,   2.699,   2.699,
  2.472,   2.472,   2.472,   2.472,
  2.788,   2.788,   2.788,   2.788,
  2.717,   2.717,   2.717,   2.717,
  2.65,    2.65,    2.65,    2.65,
  2.658,   2.658,   2.658,   2.658,
  2.913,   2.913,   2.913,   2.913,
  2.951,   2.951,   2.951,   2.951,
  2.758,   2.758,   2.758,   2.758,
  3.027,   3.027,   3.027,   3.027,
  3.261,   3.261,   3.261,   3.261,
  3.397,   3.397,   3.397,   3.397,
  3.241,   3.241,   3.241,   3.241,
  3.291,   3.291,   3.291,   3.291,
  2.969,   2.969,   2.969,   2.969,
  2.818,   2.818,   2.818,   2.818,
  2.595,   2.595,   2.595,   2.595,
  2.324,   2.324,   2.324,   2.324,
  2.327,   2.327,   2.327,   2.327,
  2.148,   2.148,   2.148,   2.148,
  2.04,    2.04,    2.04,    2.04,
  2.22,    2.22,    2.22,    2.22,
  2.112,   2.112,   2.112,   2.112,
  1.974,   1.974,   1.974,   1.974,
  2.04,    2.04,    2.04,    2.04,
  1.902,   1.902,   1.902,   1.902,
  1.937,   1.937,   1.937,   1.937,
  1.982,   1.982,   1.982,   1.982,
  2.096,   2.096,   2.096,   2.096,
  2.008,   2.008,   2.008,   2.008,
  2.02,    2.02,    2.02,    2.02,
  1.989,   1.989,   1.989,   1.989,
  1.891,   1.891,   1.891,   1.891,
  1.921,   1.921,   1.921,   1.921,
  1.884,   1.884,   1.884,   1.884,
  1.834,   1.834,   1.834,   1.834,
  1.925,   1.925,   1.925,   1.925,
  1.809,   1.809,   1.809,   1.809,
  1.685,   1.685,   1.685,   1.685,
  1.535,   1.535,   1.535,   1.535,
  1.555,   1.555,   1.555,   1.555,
  1.534,   1.534,   1.534,   1.534,
  1.805,   1.805,   1.805,   1.805,
  2.165,   2.165,   2.165,   2.165,
  2.55,    2.55,    2.55,    2.55,
  4.06,    4.06,    4.06,    4.06,
  3.91,    3.91,    3.91,    3.91,
  4.22,    4.22,    4.22,    4.22,
  3.9,     3.9,     3.9,     3.9,
  4.19,    4.19,    4.19,    4.19,
  3.98,    3.98,    3.98,    3.98,
  3.75,    3.75,    3.75,    3.75,
  3.44,    3.44,    3.44,    3.44,
  4.61,    4.61,    4.61,    4.61,
  2.913,   2.913,   2.913,   2.913,
  4.24,    4.24,    4.24,    4.24,
  4.04,    4.04,    4.04,    4.04,
  4.74,    4.74,    4.74,    4.74,
  4.61,    4.61,    4.61,    4.61,
  4.47,    4.47,    4.47,    4.47,
  4.23,    4.23,    4.23,    4.23,
  3.58,    3.58,    3.58,    3.58,
  3.9,     3.9,     3.9,     3.9,
  4.34,    4.34,    4.34,    4.34,
  3.92,    3.92,    3.92,    3.92,
  2.64,    2.64,    2.64,    2.64,
  2.57,    2.57,    2.57,    2.57,
  2.42,    2.42,    2.42,    2.42,
  1.73,    1.73,    1.73,    1.73,
  1.99,    1.99,    1.99,    1.99,
  1.88,    1.88,    1.88,    1.88,
  1.75,    1.75,    1.75,    1.75,
  1.97,    1.97,    1.97,    1.97,
  1.8,     1.8,     1.8,     1.8,
  1.21,    1.21,    1.21,    1.21,
  1.81,    1.81,    1.81,    1.81,
  1.79,    1.79,    1.79,    1.79,
  1.58,    1.58,    1.58,    1.58,
  1.41,    1.41,    1.41,    1.41,
  1.32,    1.32,    1.32,    1.32,
  1.18,    1.18,    1.18,    1.18,
  1.89,    1.89,    1.89,    1.89,
  1.83,    1.83,    1.83,    1.83,
  1.34,    1.34,    1.34,    1.34,
  1.57,    1.57,    1.57,    1.57,
  1.99,    1.99,    1.99,    1.99,
  1.35,    1.35,    1.35,    1.35,
  1.34,    1.34,    1.34,    1.34,
  1.25,    1.25,    1.25,    1.25,
  1.2,     1.2,     1.2,     1.2,
  1.27,    1.27,    1.27,    1.27,
  1.28,    1.28,    1.28,    1.28,
  1.31,    1.31,    1.31,    1.31,
  2.06,    2.06,    2.06,    2.06,
  2.03,    2.03,    2.03,    2.03,
  1.86,    1.86,    1.86,    1.86,
  2.01,    2.01,    2.01,    2.01,
  1.4,     1.4,     1.4,     1.4,
  2.34,    2.34,    2.34,    2.34,
  1.67,    1.67,    1.67,    1.67,
  1.64,    1.64,    1.64,    1.64,
  2.39,    2.39,    2.39,    2.39,
  2.8,     2.8,     2.8,     2.8,
  2.15,    2.15,    2.15,    2.15,
  1.96,    1.96,    1.96,    1.96,
  1.74,    1.74,    1.74,    1.74,
  2.91,    2.91,    2.91,    2.91,
  2.92,    2.92,    2.92,    2.92,
  2.9,     2.9,     2.9,     2.9,
  2.8,     2.8,     2.8,     2.8,
  3.25,    3.25,    3.25,    3.25,
  3.16,    3.16,    3.16,    3.16,
  2.47,    2.47,    2.47,    2.47,
  2.2,     2.2,     2.2,     2.2,
  1.97,    1.97,    1.97,    1.97,
  1.68,    1.68,    1.68,    1.68,
  1.48,    1.48,    1.48,    1.48,
  1.54,    1.54,    1.54,    1.54,
  1.6,     1.6,     1.6,     1.6,
  1.58,    1.58,    1.58,    1.58,
  1.99,    1.99,    1.99,    1.99,
  2.38,    2.38,    2.38,    2.38,
  2.34,    2.34,    2.34,    2.34,
  2.26,    2.26,    2.26,    2.26,
  2.53,    2.53,    2.53,    2.53,
  2.5,     2.5,     2.5,     2.5,
  2.48,    2.48,    2.48,    2.48,
  2.67,    2.67,    2.67,    2.67,
  2.73,    2.73,    2.73,    2.73,
  2.65,    2.65,    2.65,    2.65,
  2.72,    2.72,    2.72,    2.72,
  2.65,    2.65,    2.65,    2.65,
  2.39,    2.39,    2.39,    2.39,
  2.4,     2.4,     2.4,     2.4,
  1.95,    1.95,    1.95,    1.95,
  1.64,    1.64,    1.64,    1.64,
  1.53,    1.53,    1.53,    1.53,
  1.22,    1.22,    1.22,    1.22,
  1.05,    1.05,    1.05,    1.05,
  1.39,    1.39,    1.39,    1.39,
  1.43,    1.43,    1.43,    1.43,
  2.22,    2.22,    2.22,    2.22,
  2.08,    2.08,    2.08,    2.08,
  2.3,     2.3,     2.3,     2.3,
  2.65,    2.65,    2.65,    2.65,
  2.34,    2.34,    2.34,    2.34,
  3,       3,       3,       3,
  2.85,    2.85,    2.85,    2.85,
  2.6,     2.6,     2.6,     2.6,
  2.72,    2.72,    2.72,    2.72,
  2.72,    2.72,    2.72,    2.72,
  3.07,    3.07,    3.07,    3.07,
  2.7,     2.7,     2.7,     2.7,
  3.32,    3.32,    3.32,    3.32,
  3.41,    3.41,    3.41,    3.41,
  4.13,    4.13,    4.13,    4.13,
  3.81,    3.81,    3.81,    3.81,
  4.22,    4.22,    4.22,    4.22,
  3.65,    3.65,    3.65,    3.65,
  2.94,    2.94,    2.94,    2.94,
  3.17,    3.17,    3.17,    3.17,
  3.03,    3.03,    3.03,    3.03,
  2.55,    2.55,    2.55,    2.55,
  2.34,    2.34,    2.34,    2.34,
  2,       2,       2,       2,
  1.86,    1.86,    1.86,    1.86,
  1.69,    1.69,    1.69,    1.69,
  1.43,    1.43,    1.43,    1.43,
  1.89,    1.89,    1.89,    1.89,
  2.17,    2.17,    2.17,    2.17,
  1.78,    1.78,    1.78,    1.78,
  1.89,    1.89,    1.89,    1.89,
  2.26,    2.26,    2.26,    2.26,
  1.98,    1.98,    1.98,    1.98,
  1.7,     1.7,     1.7,     1.7,
  0.55,    0.55,    0.55,    0.55,
  0.15,    0.15,    0.15,    0.15,
  0.28,    0.28,    0.28,    0.28,
  0.37,    0.37,    0.37,    0.37,
  0.3,     0.3,     0.3,     0.3,
  0.97,    0.97,    0.97,    0.97,
  0.91,    0.91,    0.91,    0.91,
  0.86,    0.86,    0.86,    0.86,
  0.45,    0.45,    0.45,    0.45,
  1.25,    1.25,    1.25,    1.25,
  1,       1,       1,       1,
  1.11,    1.11,    1.11,    1.11,
  2.16,    2.16,    2.16,    2.16,
  2.46,    2.46,    2.46,    2.46,
  2.54,    2.54,    2.54,    2.54,
  2.54,    2.54,    2.54,    2.54,
  2.62,    2.62,    2.62,    2.62,
  2.57,    2.57,    2.57,    2.57,
  2.49,    2.49,    2.49,    2.49,
  2.52,    2.52,    2.52,    2.52,
  2.81,    2.81,    2.81,    2.81,
  3.07,    3.07,    3.07,    3.07,
  2.63,    2.63,    2.63,    2.63,
  3.11,    3.11,    3.11,    3.11,
  3.02,    3.02,    3.02,    3.02,
  3.01,    3.01,    3.01,    3.01,
  3.03,    3.03,    3.03,    3.03,
  2.49,    2.49,    2.49,    2.49,
  4.01,    4.01,    4.01,    4.01,
  4.23,    4.23,    4.23,    4.23,
  3.04,    3.04,    3.04,    3.04,
  2.78,    2.78,    2.78,    2.78,
  3.29,    3.29,    3.29,    3.29,
  2.99,    2.99,    2.99,    2.99,
  2.22,    2.22,    2.22,    2.22,
  2.28,    2.28,    2.28,    2.28,
  2.06,    2.06,    2.06,    2.06,
  1.86,    1.86,    1.86,    1.86,
  1.9,     1.9,     1.9,     1.9,
  1.94,    1.94,    1.94,    1.94,
  2,       2,       2,       2,
  2.63,    2.63,    2.63,    2.63,
  2.21,    2.21,    2.21,    2.21,
  2.37,    2.37,    2.37,    2.37,
  2.04,    2.04,    2.04,    2.04,
  1.78,    1.78,    1.78,    1.78,
  1.39,    1.39,    1.39,    1.39,
  2.33,    2.33,    2.33,    2.33,
  2.72,    2.72,    2.72,    2.72,
  2.4,     2.4,     2.4,     2.4,
  2.34,    2.34,    2.34,    2.34,
  2.22,    2.22,    2.22,    2.22,
  1.86,    1.86,    1.86,    1.86,
  1.99,    1.99,    1.99,    1.99,
  1.94,    1.94,    1.94,    1.94,
  1.45,    1.45,    1.45,    1.45,
  1.59,    1.59,    1.59,    1.59,
  2.02,    2.02,    2.02,    2.02,
  2.3,     2.3,     2.3,     2.3,
  3.58,    3.58,    3.58,    3.58,
  3.21,    3.21,    3.21,    3.21,
  3.74,    3.74,    3.74,    3.74,
  2.98,    2.98,    2.98,    2.98,
  2.76,    2.76,    2.76,    2.76,
  3.15,    3.15,    3.15,    3.15,
  3.49,    3.49,    3.49,    3.49,
  2.73,    2.73,    2.73,    2.73,
  3.93,    3.93,    3.93,    3.93,
  2.95,    2.95,    2.95,    2.95,
  2.98,    2.98,    2.98,    2.98,
  2.27,    2.27,    2.27,    2.27,
  3.29,    3.29,    3.29,    3.29,
  2.63,    2.63,    2.63,    2.63,
  2.99,    2.99,    2.99,    2.99,
  3.57,    3.57,    3.57,    3.57,
  3.83,    3.83,    3.83,    3.83,
  3.74,    3.74,    3.74,    3.74,
  3.4,     3.4,     3.4,     3.4,
  3.89,    3.89,    3.89,    3.89,
  3.14,    3.14,    3.14,    3.14,
  2.94,    2.94,    2.94,    2.94,
  2.93,    2.93,    2.93,    2.93,
  2.87,    2.87,    2.87,    2.87,
  3.28,    3.28,    3.28,    3.28,
  3.52,    3.52,    3.52,    3.52,
  3.26,    3.26,    3.26,    3.26,
  3.99,    3.99,    3.99,    3.99,
  3.62,    3.62,    3.62,    3.62,
  3.14,    3.14,    3.14,    3.14,
  2.56,    2.56,    2.56,    2.56,
  2.23,    2.23,    2.23,    2.23,
  2.17,    2.17,    2.17,    2.17,
  2.23,    2.23,    2.23,    2.23,
  2.04,    2.04,    2.04,    2.04,
  2.26,    2.26,    2.26,    2.26,
  2.1,     2.1,     2.1,     2.1,
  1.95,    1.95,    1.95,    1.95,
  2.17,    2.17,    2.17,    2.17,
  2.17,    2.17,    2.17,    2.17,
  2.25,    2.25,    2.25,    2.25,
  2.19,    2.19,    2.19,    2.19,
  2.01,    2.01,    2.01,    2.01,
  1.97,    1.97,    1.97,    1.97,
  1.79,    1.79,    1.79,    1.79,
  1.67,    1.67,    1.67,    1.67,
  1.37,    1.37,    1.37,    1.37,
  2.2,     2.2,     2.2,     2.2,
  3.19,    3.19,    3.19,    3.19,
  3.67,    3.67,    3.67,    3.67,
  4.1,     4.1,     4.1,     4.1,
  3.7,     3.7,     3.7,     3.7,
  4.43,    4.43,    4.43,    4.43,
  4.41,    4.41,    4.41,    4.41,
  4.32,    4.32,    4.32,    4.32,
  4.32,    4.32,    4.32,    4.32,
  4.55,    4.55,    4.55,    4.55,
  4.47,    4.47,    4.47,    4.47,
  3.59,    3.59,    3.59,    3.59,
  2.91,    2.91,    2.91,    2.91,
  3.18,    3.18,    3.18,    3.18,
  3.23,    3.23,    3.23,    3.23,
  2.44,    2.44,    2.44,    2.44,
  2.79,    2.79,    2.79,    2.79,
  3.6,     3.6,     3.6,     3.6,
  2.75,    2.75,    2.75,    2.75,
  2.32,    2.32,    2.32,    2.32,
  2.94,    2.94,    2.94,    2.94,
  2.3,     2.3,     2.3,     2.3,
  2.14,    2.14,    2.14,    2.14,
  1.9,     1.9,     1.9,     1.9,
  2.02,    2.02,    2.02,    2.02,
  2.43,    2.43,    2.43,    2.43,
  2.48,    2.48,    2.48,    2.48,
  2.48,    2.48,    2.48,    2.48,
  2.5,     2.5,     2.5,     2.5,
  2.5,     2.5,     2.5,     2.5,
  2.41,    2.41,    2.41,    2.41,
  2.48,    2.48,    2.48,    2.48,
  2.5,     2.5,     2.5,     2.5,
  2.26,    2.26,    2.26,    2.26,
  2.38,    2.38,    2.38,    2.38,
  2.33,    2.33,    2.33,    2.33,
  2.24,    2.24,    2.24,    2.24,
  2.36,    2.36,    2.36,    2.36,
  2.65,    2.65,    2.65,    2.65,
  2.69,    2.69,    2.69,    2.69,
  2.11,    2.11,    2.11,    2.11,
  2.08,    2.08,    2.08,    2.08,
  2.44,    2.44,    2.44,    2.44,
  2.55,    2.55,    2.55,    2.55,
  1.86,    1.86,    1.86,    1.86,
  1.44,    1.44,    1.44,    1.44,
  0.99,    0.99,    0.99,    0.99,
  0.74,    0.74,    0.74,    0.74,
  1.38,    1.38,    1.38,    1.38,
  1.2,     1.2,     1.2,     1.2,
  1.65,    1.65,    1.65,    1.65,
  1.98,    1.98,    1.98,    1.98,
  2.59,    2.59,    2.59,    2.59,
  1.96,    1.96,    1.96,    1.96,
  2.44,    2.44,    2.44,    2.44,
  2.64,    2.64,    2.64,    2.64,
  1.99,    1.99,    1.99,    1.99,
  2.14,    2.14,    2.14,    2.14,
  2.18,    2.18,    2.18,    2.18,
  2.12,    2.12,    2.12,    2.12,
  2.87,    2.87,    2.87,    2.87,
  3.28,    3.28,    3.28,    3.28,
  3.21,    3.21,    3.21,    3.21,
  2.85,    2.85,    2.85,    2.85,
  3.43,    3.43,    3.43,    3.43,
  3.21,    3.21,    3.21,    3.21,
  3.41,    3.41,    3.41,    3.41,
  3.06,    3.06,    3.06,    3.06,
  3.12,    3.12,    3.12,    3.12,
  3.3,     3.3,     3.3,     3.3,
  2.74,    2.74,    2.74,    2.74,
  2.01,    2.01,    2.01,    2.01,
  1.59,    1.59,    1.59,    1.59,
  1.66,    1.66,    1.66,    1.66,
  1.3,     1.3,     1.3,     1.3,
  1.74,    1.74,    1.74,    1.74,
  2.01,    2.01,    2.01,    2.01,
  1.92,    1.92,    1.92,    1.92,
  1.02,    1.02,    1.02,    1.02,
  1.08,    1.08,    1.08,    1.08,
  1.25,    1.25,    1.25,    1.25,
  1.74,    1.74,    1.74,    1.74,
  1.87,    1.87,    1.87,    1.87,
  1.68,    1.68,    1.68,    1.68,
  1.47,    1.47,    1.47,    1.47,
  1.74,    1.74,    1.74,    1.74,
  2.23,    2.23,    2.23,    2.23,
  1.8,     1.8,     1.8,     1.8,
  2.13,    2.13,    2.13,    2.13,
  1.66,    1.66,    1.66,    1.66,
  1.51,    1.51,    1.51,    1.51,
  1.39,    1.39,    1.39,    1.39,
  1.36,    1.36,    1.36,    1.36,
  1.84,    1.84,    1.84,    1.84,
  1.84,    1.84,    1.84,    1.84,
  1.67,    1.67,    1.67,    1.67,
  0.93,    0.93,    0.93,    0.93,
  0.97,    0.97,    0.97,    0.97,
  1.64,    1.64,    1.64,    1.64,
  2.42,    2.42,    2.42,    2.42,
  2.33,    2.33,    2.33,    2.33,
  2.38,    2.38,    2.38,    2.38,
  2.36,    2.36,    2.36,    2.36,
  2.88,    2.88,    2.88,    2.88,
  2.55,    2.55,    2.55,    2.55,
  2.44,    2.44,    2.44,    2.44,
  2.69,    2.69,    2.69,    2.69,
  2.45,    2.45,    2.45,    2.45,
  1.59,    1.59,    1.59,    1.59,
  2.89,    2.89,    2.89,    2.89,
  3.19,    3.19,    3.19,    3.19,
  2.96,    2.96,    2.96,    2.96,
  3.13,    3.13,    3.13,    3.13,
  4.45,    4.45,    4.45,    4.45,
  3.65,    3.65,    3.65,    3.65,
  3.11,    3.11,    3.11,    3.11,
  3.2,     3.2,     3.2,     3.2,
  2.49,    2.49,    2.49,    2.49,
  2.37,    2.37,    2.37,    2.37,
  2.27,    2.27,    2.27,    2.27,
  2.59,    2.59,    2.59,    2.59,
  2.13,    2.13,    2.13,    2.13,
  1.83,    1.83,    1.83,    1.83,
  1.83,    1.83,    1.83,    1.83,
  2.19,    2.19,    2.19,    2.19,
  1.89,    1.89,    1.89,    1.89,
  1.92,    1.92,    1.92,    1.92,
  1.73,    1.73,    1.73,    1.73,
  1.44,    1.44,    1.44,    1.44,
  0.76,    0.76,    0.76,    0.76,
  0.21,    0.21,    0.21,    0.21,
  0.6,     0.6,     0.6,     0.6,
  1.03,    1.03,    1.03,    1.03,
  1.71,    1.71,    1.71,    1.71,
  1.98,    1.98,    1.98,    1.98,
  1.17,    1.17,    1.17,    1.17,
  1.56,    1.56,    1.56,    1.56,
  1.42,    1.42,    1.42,    1.42,
  1.05,    1.05,    1.05,    1.05,
  1.13,    1.13,    1.13,    1.13,
  1.78,    1.78,    1.78,    1.78,
  2.08,    2.08,    2.08,    2.08,
  1.39,    1.39,    1.39,    1.39,
  1.06,    1.06,    1.06,    1.06,
  1.19,    1.19,    1.19,    1.19,
  1.65,    1.65,    1.65,    1.65,
  2.38,    2.38,    2.38,    2.38,
  2.73,    2.73,    2.73,    2.73,
  2.21,    2.21,    2.21,    2.21,
  2.94,    2.94,    2.94,    2.94,
  3.06,    3.06,    3.06,    3.06,
  2.79,    2.79,    2.79,    2.79,
  3.008,   3.008,   3.008,   3.008,
  3.267,   3.267,   3.267,   3.267,
  3.397,   3.397,   3.397,   3.397,
  3.363,   3.363,   3.363,   3.363,
  3.304,   3.304,   3.304,   3.304,
  3.289,   3.289,   3.289,   3.289,
  3.391,   3.391,   3.391,   3.391,
  3.1,     3.1,     3.1,     3.1,
  3.15,    3.15,    3.15,    3.15,
  3.36,    3.36,    3.36,    3.36,
  2.35,    2.35,    2.35,    2.35,
  2.96,    2.96,    2.96,    2.96,
  3.44,    3.44,    3.44,    3.44,
  3.39,    3.39,    3.39,    3.39,
  2.74,    2.74,    2.74,    2.74,
  2.07,    2.07,    2.07,    2.07,
  1.93,    1.93,    1.93,    1.93,
  2.21,    2.21,    2.21,    2.21,
  2.39,    2.39,    2.39,    2.39,
  2.42,    2.42,    2.42,    2.42,
  2.46,    2.46,    2.46,    2.46,
  2.35,    2.35,    2.35,    2.35,
  2.3,     2.3,     2.3,     2.3,
  1.83,    1.83,    1.83,    1.83,
  2.01,    2.01,    2.01,    2.01,
  2.54,    2.54,    2.54,    2.54,
  2.54,    2.54,    2.54,    2.54,
  2.57,    2.57,    2.57,    2.57,
  2.53,    2.53,    2.53,    2.53,
  2.58,    2.58,    2.58,    2.58,
  2.45,    2.45,    2.45,    2.45,
  2.91,    2.91,    2.91,    2.91,
  3.07,    3.07,    3.07,    3.07,
  3.02,    3.02,    3.02,    3.02,
  2.92,    2.92,    2.92,    2.92,
  2.69,    2.69,    2.69,    2.69,
  2.76,    2.76,    2.76,    2.76,
  2.99,    2.99,    2.99,    2.99,
  3.35,    3.35,    3.35,    3.35,
  3.62,    3.62,    3.62,    3.62,
  3.52,    3.52,    3.52,    3.52,
  4.61,    4.61,    4.61,    4.61,
  5,       5,       5,       5,
  4.52,    4.52,    4.52,    4.52,
  4.36,    4.36,    4.36,    4.36,
  4.91,    4.91,    4.91,    4.91,
  5.3,     5.3,     5.3,     5.3,
  4.92,    4.92,    4.92,    4.92,
  6.05,    6.05,    6.05,    6.05,
  6.18,    6.18,    6.18,    6.18,
  6.99,    6.99,    6.99,    6.99,
  6.95,    6.95,    6.95,    6.95,
  7.11,    7.11,    7.11,    7.11,
  6.85,    6.85,    6.85,    6.85,
  6.57,    6.57,    6.57,    6.57,
  6.23,    6.23,    6.23,    6.23,
  6.17,    6.17,    6.17,    6.17,
  5.77,    5.77,    5.77,    5.77,
  5.99,    5.99,    5.99,    5.99,
  6.04,    6.04,    6.04,    6.04,
  4.76,    4.76,    4.76,    4.76,
  5.16,    5.16,    5.16,    5.16,
  4.36,    4.36,    4.36,    4.36,
  3.47,    3.47,    3.47,    3.47,
  3.33,    3.33,    3.33,    3.33,
  3.2,     3.2,     3.2,     3.2,
  2.93,    2.93,    2.93,    2.93,
  3.04,    3.04,    3.04,    3.04,
  2.69,    2.69,    2.69,    2.69,
  2.69,    2.69,    2.69,    2.69,
  2.8,     2.8,     2.8,     2.8,
  2.34,    2.34,    2.34,    2.34,
  2.42,    2.42,    2.42,    2.42,
  2.35,    2.35,    2.35,    2.35,
  2.92,    2.92,    2.92,    2.92,
  2.34,    2.34,    2.34,    2.34,
  2.32,    2.32,    2.32,    2.32,
  2.02,    2.02,    2.02,    2.02,
  2,       2,       2,       2,
  1.85,    1.85,    1.85,    1.85,
  1.77,    1.77,    1.77,    1.77,
  1.58,    1.58,    1.58,    1.58,
  1.84,    1.84,    1.84,    1.84,
  1.82,    1.82,    1.82,    1.82,
  1.64,    1.64,    1.64,    1.64,
  1.74,    1.74,    1.74,    1.74,
  1.51,    1.51,    1.51,    1.51,
  1.55,    1.55,    1.55,    1.55,
  1.48,    1.48,    1.48,    1.48,
  1.43,    1.43,    1.43,    1.43,
  1.81,    1.81,    1.81,    1.81,
  1.67,    1.67,    1.67,    1.67,
  0.96,    0.96,    0.96,    0.96,
  1.18,    1.18,    1.18,    1.18,
  1.17,    1.17,    1.17,    1.17,
  1.42,    1.42,    1.42,    1.42,
  1.21,    1.21,    1.21,    1.21,
  1.39,    1.39,    1.39,    1.39,
  1.52,    1.52,    1.52,    1.52,
  1.7,     1.7,     1.7,     1.7,
  1.43,    1.43,    1.43,    1.43,
  0.03,    0.03,    0.03,    0.03,
  2.06,    2.06,    2.06,    2.06,
  2.72,    2.72,    2.72,    2.72,
  2.32,    2.32,    2.32,    2.32,
  2.59,    2.59,    2.59,    2.59,
  2.72,    2.72,    2.72,    2.72,
  2.57,    2.57,    2.57,    2.57,
  2.23,    2.23,    2.23,    2.23,
  2.6,     2.6,     2.6,     2.6,
  2.63,    2.63,    2.63,    2.63,
  2.52,    2.52,    2.52,    2.52,
  3.06,    3.06,    3.06,    3.06,
  3.14,    3.14,    3.14,    3.14,
  2.04,    2.04,    2.04,    2.04,
  1.11,    1.11,    1.11,    1.11,
  1.51,    1.51,    1.51,    1.51,
  1.67,    1.67,    1.67,    1.67,
  1.67,    1.67,    1.67,    1.67,
  2.01,    2.01,    2.01,    2.01,
  1.89,    1.89,    1.89,    1.89,
  1.89,    1.89,    1.89,    1.89,
  1.95,    1.95,    1.95,    1.95,
  2.06,    2.06,    2.06,    2.06,
  2.23,    2.23,    2.23,    2.23,
  2.38,    2.38,    2.38,    2.38,
  2.31,    2.31,    2.31,    2.31,
  2.4,     2.4,     2.4,     2.4,
  2.32,    2.32,    2.32,    2.32,
  2.29,    2.29,    2.29,    2.29,
  2.16,    2.16,    2.16,    2.16,
  2.16,    2.16,    2.16,    2.16,
  1.94,    1.94,    1.94,    1.94,
  1.91,    1.91,    1.91,    1.91,
  1.68,    1.68,    1.68,    1.68,
  1.38,    1.38,    1.38,    1.38,
  1.49,    1.49,    1.49,    1.49,
  1.91,    1.91,    1.91,    1.91,
  2.01,    2.01,    2.01,    2.01,
  2.17,    2.17,    2.17,    2.17,
  1.52,    1.52,    1.52,    1.52,
  1.24,    1.24,    1.24,    1.24,
  1.75,    1.75,    1.75,    1.75,
  2.68,    2.68,    2.68,    2.68,
  2.55,    2.55,    2.55,    2.55,
  2.61,    2.61,    2.61,    2.61,
  3.07,    3.07,    3.07,    3.07,
  2.54,    2.54,    2.54,    2.54,
  3.13,    3.13,    3.13,    3.13,
  3.36,    3.36,    3.36,    3.36,
  3.02,    3.02,    3.02,    3.02,
  3.02,    3.02,    3.02,    3.02,
  2.82,    2.82,    2.82,    2.82,
  2.12,    2.12,    2.12,    2.12,
  3.44,    3.44,    3.44,    3.44,
  2.64,    2.64,    2.64,    2.64,
  3.01,    3.01,    3.01,    3.01,
  2.38,    2.38,    2.38,    2.38,
  2.15,    2.15,    2.15,    2.15,
  2.02,    2.02,    2.02,    2.02,
  1.8,     1.8,     1.8,     1.8,
  2.06,    2.06,    2.06,    2.06,
  2.34,    2.34,    2.34,    2.34,
  1.73,    1.73,    1.73,    1.73,
  2.16,    2.16,    2.16,    2.16,
  2.63,    2.63,    2.63,    2.63,
  2.38,    2.38,    2.38,    2.38,
  2.42,    2.42,    2.42,    2.42,
  2.52,    2.52,    2.52,    2.52,
  2.29,    2.29,    2.29,    2.29,
  2.3,     2.3,     2.3,     2.3,
  2.18,    2.18,    2.18,    2.18,
  2.49,    2.49,    2.49,    2.49,
  1.93,    1.93,    1.93,    1.93,
  1.96,    1.96,    1.96,    1.96,
  2.24,    2.24,    2.24,    2.24,
  2.35,    2.35,    2.35,    2.35,
  2.45,    2.45,    2.45,    2.45,
  2.35,    2.35,    2.35,    2.35,
  2.21,    2.21,    2.21,    2.21,
  2.58,    2.58,    2.58,    2.58,
  2.36,    2.36,    2.36,    2.36,
  2.52,    2.52,    2.52,    2.52,
  2.74,    2.74,    2.74,    2.74,
  2.13,    2.13,    2.13,    2.13,
  2.69,    2.69,    2.69,    2.69,
  2.34,    2.34,    2.34,    2.34,
  1.86,    1.86,    1.86,    1.86,
  1.62,    1.62,    1.62,    1.62,
  1.71,    1.71,    1.71,    1.71,
  1.73,    1.73,    1.73,    1.73,
  1.61,    1.61,    1.61,    1.61,
  0.95,    0.95,    0.95,    0.95,
  0.47,    0.47,    0.47,    0.47,
  0.82,    0.82,    0.82,    0.82,
  0.42,    0.42,    0.42,    0.42,
  1.86,    1.86,    1.86,    1.86,
  1.69,    1.69,    1.69,    1.69,
  2.31,    2.31,    2.31,    2.31,
  2.44,    2.44,    2.44,    2.44,
  1.46,    1.46,    1.46,    1.46,
  0.94,    0.94,    0.94,    0.94,
  0.95,    0.95,    0.95,    0.95,
  0.51,    0.51,    0.51,    0.51,
  0.32,    0.32,    0.32,    0.32,
  1.14,    1.14,    1.14,    1.14,
  1.79,    1.79,    1.79,    1.79,
  1.5,     1.5,     1.5,     1.5,
  1.92,    1.92,    1.92,    1.92,
  2.24,    2.24,    2.24,    2.24,
  1.45,    1.45,    1.45,    1.45,
  1.78,    1.78,    1.78,    1.78,
  1.46,    1.46,    1.46,    1.46,
  1.56,    1.56,    1.56,    1.56,
  1.95,    1.95,    1.95,    1.95,
  2.07,    2.07,    2.07,    2.07,
  1.95,    1.95,    1.95,    1.95,
  1.98,    1.98,    1.98,    1.98,
  2.17,    2.17,    2.17,    2.17,
  2.35,    2.35,    2.35,    2.35,
  2.25,    2.25,    2.25,    2.25,
  2.51,    2.51,    2.51,    2.51,
  2.1,     2.1,     2.1,     2.1,
  2.32,    2.32,    2.32,    2.32,
  2.57,    2.57,    2.57,    2.57,
  2.54,    2.54,    2.54,    2.54,
  3.03,    3.03,    3.03,    3.03,
  2.48,    2.48,    2.48,    2.48,
  2.64,    2.64,    2.64,    2.64,
  2.87,    2.87,    2.87,    2.87,
  2.94,    2.94,    2.94,    2.94,
  3.58,    3.58,    3.58,    3.58,
  3.6,     3.6,     3.6,     3.6,
  3.13,    3.13,    3.13,    3.13,
  3.82,    3.82,    3.82,    3.82,
  3.87,    3.87,    3.87,    3.87,
  4.19,    4.19,    4.19,    4.19,
  4.03,    4.03,    4.03,    4.03,
  3.92,    3.92,    3.92,    3.92,
  4.35,    4.35,    4.35,    4.35,
  3.008,   3.008,   3.008,   3.008,
  4.47,    4.47,    4.47,    4.47,
  4.42,    4.42,    4.42,    4.42,
  4.83,    4.83,    4.83,    4.83,
  4.04,    4.04,    4.04,    4.04,
  4.45,    4.45,    4.45,    4.45,
  4.7,     4.7,     4.7,     4.7,
  4.95,    4.95,    4.95,    4.95,
  4.06,    4.06,    4.06,    4.06,
  3.93,    3.93,    3.93,    3.93,
  4.57,    4.57,    4.57,    4.57,
  5.54,    5.54,    5.54,    5.54,
  5.76,    5.76,    5.76,    5.76,
  6.01,    6.01,    6.01,    6.01,
  5.25,    5.25,    5.25,    5.25,
  5.91,    5.91,    5.91,    5.91,
  4.16,    4.16,    4.16,    4.16,
  2.88,    2.88,    2.88,    2.88,
  2.67,    2.67,    2.67,    2.67,
  3.44,    3.44,    3.44,    3.44,
  3.11,    3.11,    3.11,    3.11,
  3.54,    3.54,    3.54,    3.54,
  2.9,     2.9,     2.9,     2.9,
  4.1,     4.1,     4.1,     4.1,
  3.51,    3.51,    3.51,    3.51,
  3.67,    3.67,    3.67,    3.67,
  3.89,    3.89,    3.89,    3.89,
  4.48,    4.48,    4.48,    4.48,
  4.7,     4.7,     4.7,     4.7,
  5.18,    5.18,    5.18,    5.18,
  5.16,    5.16,    5.16,    5.16,
  4.83,    4.83,    4.83,    4.83,
  4.65,    4.65,    4.65,    4.65,
  4.26,    4.26,    4.26,    4.26,
  3.85,    3.85,    3.85,    3.85,
  3.86,    3.86,    3.86,    3.86,
  3.8,     3.8,     3.8,     3.8,
  4.08,    4.08,    4.08,    4.08,
  4.03,    4.03,    4.03,    4.03,
  4.23,    4.23,    4.23,    4.23,
  4.65,    4.65,    4.65,    4.65,
  4.79,    4.79,    4.79,    4.79,
  4.96,    4.96,    4.96,    4.96,
  4.68,    4.68,    4.68,    4.68,
  4.66,    4.66,    4.66,    4.66,
  4.9,     4.9,     4.9,     4.9,
  5.51,    5.51,    5.51,    5.51,
  5.34,    5.34,    5.34,    5.34,
  5.13,    5.13,    5.13,    5.13,
  5.4,     5.4,     5.4,     5.4,
  5.04,    5.04,    5.04,    5.04,
  5.09,    5.09,    5.09,    5.09,
  5.41,    5.41,    5.41,    5.41,
  5.46,    5.46,    5.46,    5.46,
  6.18,    6.18,    6.18,    6.18,
  5.22,    5.22,    5.22,    5.22,
  4.54,    4.54,    4.54,    4.54,
  4.69,    4.69,    4.69,    4.69,
  4.82,    4.82,    4.82,    4.82,
  4.97,    4.97,    4.97,    4.97,
  4.55,    4.55,    4.55,    4.55,
  4.85,    4.85,    4.85,    4.85,
  3.84,    3.84,    3.84,    3.84,
  4.46,    4.46,    4.46,    4.46,
  3.88,    3.88,    3.88,    3.88,
  3.87,    3.87,    3.87,    3.87,
  3.54,    3.54,    3.54,    3.54,
  3.34,    3.34,    3.34,    3.34,
  3.43,    3.43,    3.43,    3.43,
  2.85,    2.85,    2.85,    2.85,
  2.67,    2.67,    2.67,    2.67,
  3.29,    3.29,    3.29,    3.29,
  3.54,    3.54,    3.54,    3.54,
  3.16,    3.16,    3.16,    3.16,
  2.99,    2.99,    2.99,    2.99,
  3.55,    3.55,    3.55,    3.55,
  2.92,    2.92,    2.92,    2.92,
  3.18,    3.18,    3.18,    3.18,
  2.7,     2.7,     2.7,     2.7,
  2.24,    2.24,    2.24,    2.24,
  1.88,    1.88,    1.88,    1.88,
  1.72,    1.72,    1.72,    1.72,
  1.1,     1.1,     1.1,     1.1,
  1.72,    1.72,    1.72,    1.72,
  2.12,    2.12,    2.12,    2.12,
  2.47,    2.47,    2.47,    2.47,
  2.36,    2.36,    2.36,    2.36,
  2.9,     2.9,     2.9,     2.9,
  2.27,    2.27,    2.27,    2.27,
  2.42,    2.42,    2.42,    2.42,
  3.02,    3.02,    3.02,    3.02,
  2.94,    2.94,    2.94,    2.94,
  2.98,    2.98,    2.98,    2.98,
  3.32,    3.32,    3.32,    3.32,
  3.31,    3.31,    3.31,    3.31,
  3.19,    3.19,    3.19,    3.19,
  3.37,    3.37,    3.37,    3.37,
  3.26,    3.26,    3.26,    3.26,
  3.7,     3.7,     3.7,     3.7,
  3.17,    3.17,    3.17,    3.17,
  2.75,    2.75,    2.75,    2.75,
  2.88,    2.88,    2.88,    2.88,
  2.83,    2.83,    2.83,    2.83,
  3.3,     3.3,     3.3,     3.3,
  2.82,    2.82,    2.82,    2.82,
  2.87,    2.87,    2.87,    2.87,
  2.93,    2.93,    2.93,    2.93,
  2.75,    2.75,    2.75,    2.75,
  2.49,    2.49,    2.49,    2.49,
  1.7,     1.7,     1.7,     1.7,
  1.56,    1.56,    1.56,    1.56,
  1.6,     1.6,     1.6,     1.6,
  1.31,    1.31,    1.31,    1.31,
  1.23,    1.23,    1.23,    1.23,
  1.63,    1.63,    1.63,    1.63,
  1.98,    1.98,    1.98,    1.98,
  1.77,    1.77,    1.77,    1.77,
  1.96,    1.96,    1.96,    1.96,
  1.79,    1.79,    1.79,    1.79,
  1.84,    1.84,    1.84,    1.84,
  1.16,    1.16,    1.16,    1.16,
  0.62,    0.62,    0.62,    0.62,
  0.58,    0.58,    0.58,    0.58,
  0.85,    0.85,    0.85,    0.85,
  1.65,    1.65,    1.65,    1.65,
  0.6,     0.6,     0.6,     0.6,
  0.87,    0.87,    0.87,    0.87,
  0.58,    0.58,    0.58,    0.58,
  0.81,    0.81,    0.81,    0.81,
  1.12,    1.12,    1.12,    1.12,
  0.63,    0.63,    0.63,    0.63,
  1.11,    1.11,    1.11,    1.11,
  1.29,    1.29,    1.29,    1.29,
  1.16,    1.16,    1.16,    1.16,
  0.57,    0.57,    0.57,    0.57,
  0.4,     0.4,     0.4,     0.4,
  0.37,    0.37,    0.37,    0.37,
  0.57,    0.57,    0.57,    0.57,
  1.13,    1.13,    1.13,    1.13,
  1.37,    1.37,    1.37,    1.37,
  1.89,    1.89,    1.89,    1.89,
  1.19,    1.19,    1.19,    1.19,
  1.42,    1.42,    1.42,    1.42,
  2.06,    2.06,    2.06,    2.06,
  1.26,    1.26,    1.26,    1.26,
  1.2,     1.2,     1.2,     1.2,
  1.53,    1.53,    1.53,    1.53,
  2.31,    2.31,    2.31,    2.31,
  1.76,    1.76,    1.76,    1.76,
  1.9,     1.9,     1.9,     1.9,
  1.71,    1.71,    1.71,    1.71,
  1.01,    1.01,    1.01,    1.01,
  1.26,    1.26,    1.26,    1.26,
  0.86,    0.86,    0.86,    0.86,
  0.57,    0.57,    0.57,    0.57,
  0.91,    0.91,    0.91,    0.91,
  0.77,    0.77,    0.77,    0.77,
  0.28,    0.28,    0.28,    0.28,
  1.05,    1.05,    1.05,    1.05,
  0.99,    0.99,    0.99,    0.99,
  1.58,    1.58,    1.58,    1.58,
  1.86,    1.86,    1.86,    1.86,
  1.89,    1.89,    1.89,    1.89,
  1.87,    1.87,    1.87,    1.87,
  1.74,    1.74,    1.74,    1.74,
  1.15,    1.15,    1.15,    1.15,
  1.34,    1.34,    1.34,    1.34,
  1.53,    1.53,    1.53,    1.53,
  1.31,    1.31,    1.31,    1.31,
  1.22,    1.22,    1.22,    1.22,
  1.52,    1.52,    1.52,    1.52,
  1.57,    1.57,    1.57,    1.57,
  1.48,    1.48,    1.48,    1.48,
  1.31,    1.31,    1.31,    1.31,
  1.68,    1.68,    1.68,    1.68,
  2.32,    2.32,    2.32,    2.32,
  2.43,    2.43,    2.43,    2.43,
  2.26,    2.26,    2.26,    2.26,
  2.15,    2.15,    2.15,    2.15,
  1.74,    1.74,    1.74,    1.74,
  1.72,    1.72,    1.72,    1.72,
  1.64,    1.64,    1.64,    1.64,
  1.29,    1.29,    1.29,    1.29,
  1.22,    1.22,    1.22,    1.22,
  1.12,    1.12,    1.12,    1.12,
  1.78,    1.78,    1.78,    1.78,
  2.16,    2.16,    2.16,    2.16,
  2.07,    2.07,    2.07,    2.07,
  2.03,    2.03,    2.03,    2.03,
  2.42,    2.42,    2.42,    2.42,
  2.11,    2.11,    2.11,    2.11,
  2.29,    2.29,    2.29,    2.29,
  2.19,    2.19,    2.19,    2.19,
  2.45,    2.45,    2.45,    2.45,
  2.37,    2.37,    2.37,    2.37,
  2.6,     2.6,     2.6,     2.6,
  2.17,    2.17,    2.17,    2.17,
  2.05,    2.05,    2.05,    2.05,
  2.79,    2.79,    2.79,    2.79,
  2.63,    2.63,    2.63,    2.63,
  2.21,    2.21,    2.21,    2.21,
  1.97,    1.97,    1.97,    1.97,
  1.25,    1.25,    1.25,    1.25,
  2.03,    2.03,    2.03,    2.03,
  2,       2,       2,       2,
  1.84,    1.84,    1.84,    1.84,
  2.16,    2.16,    2.16,    2.16,
  1.88,    1.88,    1.88,    1.88,
  1.56,    1.56,    1.56,    1.56,
  2.06,    2.06,    2.06,    2.06,
  2.02,    2.02,    2.02,    2.02,
  1.5,     1.5,     1.5,     1.5,
  1.81,    1.81,    1.81,    1.81,
  1.33,    1.33,    1.33,    1.33,
  1.12,    1.12,    1.12,    1.12,
  1.18,    1.18,    1.18,    1.18,
  2.04,    2.04,    2.04,    2.04,
  2.57,    2.57,    2.57,    2.57,
  2.33,    2.33,    2.33,    2.33,
  0.53,    0.53,    0.53,    0.53,
  2.31,    2.31,    2.31,    2.31,
  1.9,     1.9,     1.9,     1.9,
  2.18,    2.18,    2.18,    2.18,
  1.98,    1.98,    1.98,    1.98,
  2.37,    2.37,    2.37,    2.37,
  1.8,     1.8,     1.8,     1.8,
  2.29,    2.29,    2.29,    2.29,
  2.13,    2.13,    2.13,    2.13,
  2.69,    2.69,    2.69,    2.69,
  2.89,    2.89,    2.89,    2.89,
  2.82,    2.82,    2.82,    2.82,
  1.6,     1.6,     1.6,     1.6,
  1.8,     1.8,     1.8,     1.8,
  2.33,    2.33,    2.33,    2.33,
  2.32,    2.32,    2.32,    2.32,
  2.28,    2.28,    2.28,    2.28,
  2.3,     2.3,     2.3,     2.3,
  2.05,    2.05,    2.05,    2.05,
  2.23,    2.23,    2.23,    2.23,
  1.97,    1.97,    1.97,    1.97,
  2.1,     2.1,     2.1,     2.1,
  2.07,    2.07,    2.07,    2.07,
  1.48,    1.48,    1.48,    1.48,
  1.86,    1.86,    1.86,    1.86,
  1.3,     1.3,     1.3,     1.3,
  2.01,    2.01,    2.01,    2.01,
  1.09,    1.09,    1.09,    1.09,
  1.31,    1.31,    1.31,    1.31,
  1.34,    1.34,    1.34,    1.34,
  1.67,    1.67,    1.67,    1.67,
  2.58,    2.58,    2.58,    2.58,
  3.31,    3.31,    3.31,    3.31,
  3.48,    3.48,    3.48,    3.48,
  3.42,    3.42,    3.42,    3.42,
  3.51,    3.51,    3.51,    3.51,
  3.48,    3.48,    3.48,    3.48,
  3.33,    3.33,    3.33,    3.33,
  2.66,    2.66,    2.66,    2.66,
  2.48,    2.48,    2.48,    2.48,
  2.86,    2.86,    2.86,    2.86,
  3.03,    3.03,    3.03,    3.03,
  3.01,    3.01,    3.01,    3.01,
  2.3,     2.3,     2.3,     2.3,
  2.5,     2.5,     2.5,     2.5,
  2.12,    2.12,    2.12,    2.12,
  0.73,    0.73,    0.73,    0.73,
  1.39,    1.39,    1.39,    1.39,
  1.61,    1.61,    1.61,    1.61,
  1.07,    1.07,    1.07,    1.07,
  1.34,    1.34,    1.34,    1.34,
  1.4,     1.4,     1.4,     1.4,
  1.3,     1.3,     1.3,     1.3,
  2.09,    2.09,    2.09,    2.09,
  1.85,    1.85,    1.85,    1.85,
  2.76,    2.76,    2.76,    2.76,
  2.67,    2.67,    2.67,    2.67,
  2.37,    2.37,    2.37,    2.37,
  2.19,    2.19,    2.19,    2.19,
  3.49,    3.49,    3.49,    3.49,
  3.25,    3.25,    3.25,    3.25,
  3.42,    3.42,    3.42,    3.42,
  4,       4,       4,       4,
  3.98,    3.98,    3.98,    3.98,
  3.74,    3.74,    3.74,    3.74,
  3.4,     3.4,     3.4,     3.4,
  4.42,    4.42,    4.42,    4.42,
  4.57,    4.57,    4.57,    4.57,
  4.51,    4.51,    4.51,    4.51,
  4.09,    4.09,    4.09,    4.09,
  4.9,     4.9,     4.9,     4.9,
  5.23,    5.23,    5.23,    5.23,
  4.28,    4.28,    4.28,    4.28,
  3.74,    3.74,    3.74,    3.74,
  4.62,    4.62,    4.62,    4.62,
  4.31,    4.31,    4.31,    4.31,
  3.65,    3.65,    3.65,    3.65,
  4.11,    4.11,    4.11,    4.11,
  4.21,    4.21,    4.21,    4.21,
  3.66,    3.66,    3.66,    3.66,
  3.68,    3.68,    3.68,    3.68,
  3.79,    3.79,    3.79,    3.79,
  4.1,     4.1,     4.1,     4.1,
  4.19,    4.19,    4.19,    4.19,
  4.03,    4.03,    4.03,    4.03,
  4.4,     4.4,     4.4,     4.4,
  4.62,    4.62,    4.62,    4.62,
  4.27,    4.27,    4.27,    4.27,
  3.9,     3.9,     3.9,     3.9,
  4.37,    4.37,    4.37,    4.37,
  5.02,    5.02,    5.02,    5.02,
  4.48,    4.48,    4.48,    4.48,
  3.89,    3.89,    3.89,    3.89,
  3.22,    3.22,    3.22,    3.22,
  3.16,    3.16,    3.16,    3.16,
  3.3,     3.3,     3.3,     3.3,
  2.22,    2.22,    2.22,    2.22,
  2.06,    2.06,    2.06,    2.06,
  2.32,    2.32,    2.32,    2.32,
  2.82,    2.82,    2.82,    2.82,
  2.75,    2.75,    2.75,    2.75,
  2.77,    2.77,    2.77,    2.77,
  2.1,     2.1,     2.1,     2.1,
  1.56,    1.56,    1.56,    1.56,
  1.84,    1.84,    1.84,    1.84,
  1.89,    1.89,    1.89,    1.89,
  1.79,    1.79,    1.79,    1.79,
  2.08,    2.08,    2.08,    2.08,
  1.73,    1.73,    1.73,    1.73,
  1.89,    1.89,    1.89,    1.89,
  1.97,    1.97,    1.97,    1.97,
  2.22,    2.22,    2.22,    2.22,
  1.72,    1.72,    1.72,    1.72,
  2.19,    2.19,    2.19,    2.19,
  3.23,    3.23,    3.23,    3.23,
  3.56,    3.56,    3.56,    3.56,
  3.18,    3.18,    3.18,    3.18,
  3.9,     3.9,     3.9,     3.9,
  4.16,    4.16,    4.16,    4.16,
  4.4,     4.4,     4.4,     4.4,
  4.26,    4.26,    4.26,    4.26,
  4.06,    4.06,    4.06,    4.06,
  3.18,    3.18,    3.18,    3.18,
  2.67,    2.67,    2.67,    2.67,
  2.26,    2.26,    2.26,    2.26,
  1.81,    1.81,    1.81,    1.81,
  3.11,    3.11,    3.11,    3.11,
  3.46,    3.46,    3.46,    3.46,
  3.4,     3.4,     3.4,     3.4,
  3.5,     3.5,     3.5,     3.5,
  3.35,    3.35,    3.35,    3.35,
  2.77,    2.77,    2.77,    2.77,
  2.56,    2.56,    2.56,    2.56,
  2.67,    2.67,    2.67,    2.67,
  3.12,    3.12,    3.12,    3.12,
  2.66,    2.66,    2.66,    2.66,
  2.54,    2.54,    2.54,    2.54,
  2.92,    2.92,    2.92,    2.92,
  3.07,    3.07,    3.07,    3.07,
  3.02,    3.02,    3.02,    3.02,
  3.11,    3.11,    3.11,    3.11,
  2.22,    2.22,    2.22,    2.22,
  3.05,    3.05,    3.05,    3.05,
  2.85,    2.85,    2.85,    2.85,
  3.08,    3.08,    3.08,    3.08,
  3.65,    3.65,    3.65,    3.65,
  3.96,    3.96,    3.96,    3.96,
  3.7,     3.7,     3.7,     3.7,
  3.7,     3.7,     3.7,     3.7,
  3.39,    3.39,    3.39,    3.39,
  2.9,     2.9,     2.9,     2.9,
  3.39,    3.39,    3.39,    3.39,
  3.41,    3.41,    3.41,    3.41,
  3.06,    3.06,    3.06,    3.06,
  3.72,    3.72,    3.72,    3.72,
  3.85,    3.85,    3.85,    3.85,
  3.63,    3.63,    3.63,    3.63,
  3.77,    3.77,    3.77,    3.77,
  4.2,     4.2,     4.2,     4.2,
  3.31,    3.31,    3.31,    3.31,
  3.32,    3.32,    3.32,    3.32,
  3.31,    3.31,    3.31,    3.31,
  2.96,    2.96,    2.96,    2.96,
  3.29,    3.29,    3.29,    3.29,
  2.81,    2.81,    2.81,    2.81,
  3.3,     3.3,     3.3,     3.3,
  3.91,    3.91,    3.91,    3.91,
  3.59,    3.59,    3.59,    3.59,
  3.71,    3.71,    3.71,    3.71,
  4.19,    4.19,    4.19,    4.19,
  4.28,    4.28,    4.28,    4.28,
  3.84,    3.84,    3.84,    3.84,
  3.53,    3.53,    3.53,    3.53,
  3.67,    3.67,    3.67,    3.67,
  3.14,    3.14,    3.14,    3.14,
  2.98,    2.98,    2.98,    2.98,
  2.57,    2.57,    2.57,    2.57,
  2.54,    2.54,    2.54,    2.54,
  3.3,     3.3,     3.3,     3.3,
  2.73,    2.73,    2.73,    2.73,
  2.9,     2.9,     2.9,     2.9,
  2.96,    2.96,    2.96,    2.96,
  2.76,    2.76,    2.76,    2.76,
  1.68,    1.68,    1.68,    1.68,
  1.77,    1.77,    1.77,    1.77,
  2.09,    2.09,    2.09,    2.09,
  2.32,    2.32,    2.32,    2.32,
  2.6,     2.6,     2.6,     2.6,
  2.89,    2.89,    2.89,    2.89,
  2.99,    2.99,    2.99,    2.99,
  2.22,    2.22,    2.22,    2.22,
  2.25,    2.25,    2.25,    2.25,
  2.36,    2.36,    2.36,    2.36,
  2.65,    2.65,    2.65,    2.65,
  2.69,    2.69,    2.69,    2.69,
  2.23,    2.23,    2.23,    2.23,
  0.93,    0.93,    0.93,    0.93,
  2.63,    2.63,    2.63,    2.63,
  1.99,    1.99,    1.99,    1.99,
  2.39,    2.39,    2.39,    2.39,
  2.05,    2.05,    2.05,    2.05,
  2.06,    2.06,    2.06,    2.06,
  2.04,    2.04,    2.04,    2.04,
  2.33,    2.33,    2.33,    2.33,
  2.63,    2.63,    2.63,    2.63,
  3.2,     3.2,     3.2,     3.2,
  3.49,    3.49,    3.49,    3.49,
  3.7,     3.7,     3.7,     3.7,
  4.11,    4.11,    4.11,    4.11,
  4.08,    4.08,    4.08,    4.08,
  3.45,    3.45,    3.45,    3.45,
  4.29,    4.29,    4.29,    4.29,
  1.27,    1.27,    1.27,    1.27,
  3.01,    3.01,    3.01,    3.01,
  3.23,    3.23,    3.23,    3.23,
  4.04,    4.04,    4.04,    4.04,
  3.46,    3.46,    3.46,    3.46,
  2.09,    2.09,    2.09,    2.09,
  3.38,    3.38,    3.38,    3.38,
  1.85,    1.85,    1.85,    1.85,
  2.05,    2.05,    2.05,    2.05,
  1.54,    1.54,    1.54,    1.54,
  1.46,    1.46,    1.46,    1.46,
  2.39,    2.39,    2.39,    2.39,
  2.96,    2.96,    2.96,    2.96,
  2.27,    2.27,    2.27,    2.27,
  1.38,    1.38,    1.38,    1.38,
  0.67,    0.67,    0.67,    0.67,
  0.79,    0.79,    0.79,    0.79,
  1.05,    1.05,    1.05,    1.05,
  1.76,    1.76,    1.76,    1.76,
  2.06,    2.06,    2.06,    2.06,
  2.05,    2.05,    2.05,    2.05,
  2.31,    2.31,    2.31,    2.31,
  1.87,    1.87,    1.87,    1.87,
  1.94,    1.94,    1.94,    1.94,
  2.37,    2.37,    2.37,    2.37,
  2.28,    2.28,    2.28,    2.28,
  2.16,    2.16,    2.16,    2.16,
  2.32,    2.32,    2.32,    2.32,
  2.26,    2.26,    2.26,    2.26,
  2.32,    2.32,    2.32,    2.32,
  2.44,    2.44,    2.44,    2.44,
  2.42,    2.42,    2.42,    2.42,
  2.21,    2.21,    2.21,    2.21,
  2.27,    2.27,    2.27,    2.27,
  2.37,    2.37,    2.37,    2.37,
  2.33,    2.33,    2.33,    2.33,
  2.8,     2.8,     2.8,     2.8,
  2.91,    2.91,    2.91,    2.91,
  3.45,    3.45,    3.45,    3.45,
  3.4,     3.4,     3.4,     3.4,
  3.63,    3.63,    3.63,    3.63,
  4.07,    4.07,    4.07,    4.07,
  4.98,    4.98,    4.98,    4.98,
  5.03,    5.03,    5.03,    5.03,
  5.1,     5.1,     5.1,     5.1,
  5.58,    5.58,    5.58,    5.58,
  5.47,    5.47,    5.47,    5.47,
  5.92,    5.92,    5.92,    5.92,
  5.63,    5.63,    5.63,    5.63,
  4.81,    4.81,    4.81,    4.81,
  4.17,    4.17,    4.17,    4.17,
  4.81,    4.81,    4.81,    4.81,
  4.47,    4.47,    4.47,    4.47,
  5.57,    5.57,    5.57,    5.57,
  5.01,    5.01,    5.01,    5.01,
  4.34,    4.34,    4.34,    4.34,
  4.84,    4.84,    4.84,    4.84,
  3.41,    3.41,    3.41,    3.41,
  4,       4,       4,       4,
  3.66,    3.66,    3.66,    3.66,
  2.64,    2.64,    2.64,    2.64,
  2.78,    2.78,    2.78,    2.78,
  2.39,    2.39,    2.39,    2.39,
  3.1,     3.1,     3.1,     3.1,
  2.93,    2.93,    2.93,    2.93,
  2.59,    2.59,    2.59,    2.59,
  2.7,     2.7,     2.7,     2.7,
  3.22,    3.22,    3.22,    3.22,
  2.89,    2.89,    2.89,    2.89,
  2.72,    2.72,    2.72,    2.72,
  3.08,    3.08,    3.08,    3.08,
  2.79,    2.79,    2.79,    2.79,
  2.93,    2.93,    2.93,    2.93,
  3.31,    3.31,    3.31,    3.31,
  3.57,    3.57,    3.57,    3.57,
  2.89,    2.89,    2.89,    2.89,
  3.3,     3.3,     3.3,     3.3,
  3.21,    3.21,    3.21,    3.21,
  3.32,    3.32,    3.32,    3.32,
  3.61,    3.61,    3.61,    3.61,
  3.69,    3.69,    3.69,    3.69,
  3.54,    3.54,    3.54,    3.54,
  3.59,    3.59,    3.59,    3.59,
  3.75,    3.75,    3.75,    3.75,
  3.6,     3.6,     3.6,     3.6,
  3.45,    3.45,    3.45,    3.45,
  3.26,    3.26,    3.26,    3.26,
  3.07,    3.07,    3.07,    3.07,
  2.95,    2.95,    2.95,    2.95,
  3.44,    3.44,    3.44,    3.44,
  3.57,    3.57,    3.57,    3.57,
  3.21,    3.21,    3.21,    3.21,
  2.84,    2.84,    2.84,    2.84,
  2.51,    2.51,    2.51,    2.51,
  3.41,    3.41,    3.41,    3.41,
  3.44,    3.44,    3.44,    3.44,
  2.64,    2.64,    2.64,    2.64,
  3.32,    3.32,    3.32,    3.32,
  4.23,    4.23,    4.23,    4.23,
  4.08,    4.08,    4.08,    4.08,
  4.19,    4.19,    4.19,    4.19,
  4.81,    4.81,    4.81,    4.81,
  5.52,    5.52,    5.52,    5.52,
  4.6,     4.6,     4.6,     4.6,
  5.54,    5.54,    5.54,    5.54,
  4.85,    4.85,    4.85,    4.85,
  4.48,    4.48,    4.48,    4.48,
  4.6,     4.6,     4.6,     4.6,
  3.67,    3.67,    3.67,    3.67,
  2.42,    2.42,    2.42,    2.42,
  3.82,    3.82,    3.82,    3.82,
  3.17,    3.17,    3.17,    3.17,
  2.93,    2.93,    2.93,    2.93,
  2.12,    2.12,    2.12,    2.12,
  2.46,    2.46,    2.46,    2.46,
  2.5,     2.5,     2.5,     2.5,
  2.58,    2.58,    2.58,    2.58,
  2.48,    2.48,    2.48,    2.48,
  2.39,    2.39,    2.39,    2.39,
  2.51,    2.51,    2.51,    2.51,
  2.39,    2.39,    2.39,    2.39,
  2.47,    2.47,    2.47,    2.47,
  2.71,    2.71,    2.71,    2.71,
  3.11,    3.11,    3.11,    3.11,
  2.62,    2.62,    2.62,    2.62,
  2.48,    2.48,    2.48,    2.48,
  2.57,    2.57,    2.57,    2.57,
  3.28,    3.28,    3.28,    3.28,
  3.44,    3.44,    3.44,    3.44,
  3.27,    3.27,    3.27,    3.27,
  3.58,    3.58,    3.58,    3.58,
  3.09,    3.09,    3.09,    3.09,
  3.65,    3.65,    3.65,    3.65,
  3.8,     3.8,     3.8,     3.8,
  3.33,    3.33,    3.33,    3.33,
  3.2,     3.2,     3.2,     3.2,
  3.54,    3.54,    3.54,    3.54,
  3.79,    3.79,    3.79,    3.79,
  3.66,    3.66,    3.66,    3.66,
  3.9,     3.9,     3.9,     3.9,
  4.11,    4.11,    4.11,    4.11,
  4.11,    4.11,    4.11,    4.11,
  4.02,    4.02,    4.02,    4.02,
  4.22,    4.22,    4.22,    4.22,
  4.25,    4.25,    4.25,    4.25,
  2.74,    2.74,    2.74,    2.74,
  4.46,    4.46,    4.46,    4.46,
  4.85,    4.85,    4.85,    4.85,
  4.55,    4.55,    4.55,    4.55,
  4.02,    4.02,    4.02,    4.02,
  4.45,    4.45,    4.45,    4.45,
  4.68,    4.68,    4.68,    4.68,
  4.52,    4.52,    4.52,    4.52,
  4.26,    4.26,    4.26,    4.26,
  5.02,    5.02,    5.02,    5.02,
  4.45,    4.45,    4.45,    4.45,
  4.51,    4.51,    4.51,    4.51,
  4.03,    4.03,    4.03,    4.03,
  4.46,    4.46,    4.46,    4.46,
  3.82,    3.82,    3.82,    3.82,
  4.21,    4.21,    4.21,    4.21,
  4.23,    4.23,    4.23,    4.23,
  4.25,    4.25,    4.25,    4.25,
  4.17,    4.17,    4.17,    4.17,
  4.92,    4.92,    4.92,    4.92,
  4.12,    4.12,    4.12,    4.12,
  3.5,     3.5,     3.5,     3.5,
  3.14,    3.14,    3.14,    3.14,
  3.84,    3.84,    3.84,    3.84,
  4.48,    4.48,    4.48,    4.48,
  2.94,    2.94,    2.94,    2.94,
  2.74,    2.74,    2.74,    2.74,
  3.08,    3.08,    3.08,    3.08,
  2.79,    2.79,    2.79,    2.79,
  2.5,     2.5,     2.5,     2.5,
  2.49,    2.49,    2.49,    2.49,
  1.71,    1.71,    1.71,    1.71,
  1.75,    1.75,    1.75,    1.75,
  2.12,    2.12,    2.12,    2.12,
  2.09,    2.09,    2.09,    2.09,
  2.27,    2.27,    2.27,    2.27,
  2.35,    2.35,    2.35,    2.35,
  2.72,    2.72,    2.72,    2.72,
  2.61,    2.61,    2.61,    2.61,
  3.39,    3.39,    3.39,    3.39,
  3.49,    3.49,    3.49,    3.49,
  3.91,    3.91,    3.91,    3.91,
  4.43,    4.43,    4.43,    4.43,
  4.93,    4.93,    4.93,    4.93,
  5.05,    5.05,    5.05,    5.05,
  4.68,    4.68,    4.68,    4.68,
  5.04,    5.04,    5.04,    5.04,
  4.54,    4.54,    4.54,    4.54,
  4.29,    4.29,    4.29,    4.29,
  4.35,    4.35,    4.35,    4.35,
  4.73,    4.73,    4.73,    4.73,
  5.32,    5.32,    5.32,    5.32,
  3.96,    3.96,    3.96,    3.96,
  5.04,    5.04,    5.04,    5.04,
  4.2,     4.2,     4.2,     4.2,
  3.9,     3.9,     3.9,     3.9,
  2.57,    2.57,    2.57,    2.57,
  2.01,    2.01,    2.01,    2.01,
  2.57,    2.57,    2.57,    2.57,
  3.66,    3.66,    3.66,    3.66,
  3.73,    3.73,    3.73,    3.73,
  3.77,    3.77,    3.77,    3.77,
  2.53,    2.53,    2.53,    2.53,
  2.07,    2.07,    2.07,    2.07,
  1.91,    1.91,    1.91,    1.91,
  1.92,    1.92,    1.92,    1.92,
  2.42,    2.42,    2.42,    2.42,
  2.58,    2.58,    2.58,    2.58,
  2.63,    2.63,    2.63,    2.63,
  2.74,    2.74,    2.74,    2.74,
  2.9,     2.9,     2.9,     2.9,
  2.79,    2.79,    2.79,    2.79,
  2.73,    2.73,    2.73,    2.73,
  2.2,     2.2,     2.2,     2.2,
  2.48,    2.48,    2.48,    2.48,
  2.82,    2.82,    2.82,    2.82,
  3.1,     3.1,     3.1,     3.1,
  2.99,    2.99,    2.99,    2.99,
  2.6,     2.6,     2.6,     2.6,
  2.65,    2.65,    2.65,    2.65,
  2.71,    2.71,    2.71,    2.71,
  2.95,    2.95,    2.95,    2.95,
  2.92,    2.92,    2.92,    2.92,
  3.21,    3.21,    3.21,    3.21,
  3.3,     3.3,     3.3,     3.3,
  3.42,    3.42,    3.42,    3.42,
  3.68,    3.68,    3.68,    3.68,
  3.73,    3.73,    3.73,    3.73,
  3.74,    3.74,    3.74,    3.74,
  4.47,    4.47,    4.47,    4.47,
  4.33,    4.33,    4.33,    4.33,
  4.75,    4.75,    4.75,    4.75,
  4.78,    4.78,    4.78,    4.78,
  4.76,    4.76,    4.76,    4.76,
  4.76,    4.76,    4.76,    4.76,
  4.08,    4.08,    4.08,    4.08,
  4.23,    4.23,    4.23,    4.23,
  4.2,     4.2,     4.2,     4.2,
  3.84,    3.84,    3.84,    3.84,
  4.05,    4.05,    4.05,    4.05,
  4.57,    4.57,    4.57,    4.57,
  4.64,    4.64,    4.64,    4.64,
  4.83,    4.83,    4.83,    4.83,
  3.89,    3.89,    3.89,    3.89,
  4.18,    4.18,    4.18,    4.18,
  3.55,    3.55,    3.55,    3.55,
  4.39,    4.39,    4.39,    4.39,
  4.29,    4.29,    4.29,    4.29,
  4.51,    4.51,    4.51,    4.51,
  3.98,    3.98,    3.98,    3.98,
  2.38,    2.38,    2.38,    2.38,
  1.59,    1.59,    1.59,    1.59,
  1.66,    1.66,    1.66,    1.66,
  1.73,    1.73,    1.73,    1.73,
  1.45,    1.45,    1.45,    1.45,
  1.9,     1.9,     1.9,     1.9,
  2.03,    2.03,    2.03,    2.03,
  2.22,    2.22,    2.22,    2.22,
  2.05,    2.05,    2.05,    2.05,
  2.16,    2.16,    2.16,    2.16,
  2.13,    2.13,    2.13,    2.13,
  2.27,    2.27,    2.27,    2.27,
  2.03,    2.03,    2.03,    2.03,
  2.27,    2.27,    2.27,    2.27,
  2.23,    2.23,    2.23,    2.23,
  1.96,    1.96,    1.96,    1.96,
  2.09,    2.09,    2.09,    2.09,
  2.15,    2.15,    2.15,    2.15,
  2.01,    2.01,    2.01,    2.01,
  2.13,    2.13,    2.13,    2.13,
  1.71,    1.71,    1.71,    1.71,
  1.16,    1.16,    1.16,    1.16,
  0.59,    0.59,    0.59,    0.59,
  0.85,    0.85,    0.85,    0.85,
  1.39,    1.39,    1.39,    1.39,
  1.14,    1.14,    1.14,    1.14,
  1.51,    1.51,    1.51,    1.51,
  1.66,    1.66,    1.66,    1.66,
  2.15,    2.15,    2.15,    2.15,
  1.36,    1.36,    1.36,    1.36,
  1.8,     1.8,     1.8,     1.8,
  2.53,    2.53,    2.53,    2.53,
  2.93,    2.93,    2.93,    2.93,
  3.33,    3.33,    3.33,    3.33,
  2.67,    2.67,    2.67,    2.67,
  3.62,    3.62,    3.62,    3.62,
  2.56,    2.56,    2.56,    2.56,
  3.01,    3.01,    3.01,    3.01,
  3.74,    3.74,    3.74,    3.74,
  1.9,     1.9,     1.9,     1.9,
  2.19,    2.19,    2.19,    2.19,
  2.42,    2.42,    2.42,    2.42,
  1.81,    1.81,    1.81,    1.81,
  1.95,    1.95,    1.95,    1.95,
  2.03,    2.03,    2.03,    2.03,
  2.41,    2.41,    2.41,    2.41,
  2.67,    2.67,    2.67,    2.67,
  2.91,    2.91,    2.91,    2.91,
  2.11,    2.11,    2.11,    2.11,
  1.46,    1.46,    1.46,    1.46,
  1.71,    1.71,    1.71,    1.71,
  2.01,    2.01,    2.01,    2.01,
  2.23,    2.23,    2.23,    2.23,
  2.33,    2.33,    2.33,    2.33,
  2.33,    2.33,    2.33,    2.33,
  2.37,    2.37,    2.37,    2.37,
  2.15,    2.15,    2.15,    2.15,
  2.11,    2.11,    2.11,    2.11,
  1.53,    1.53,    1.53,    1.53,
  1.93,    1.93,    1.93,    1.93,
  1.95,    1.95,    1.95,    1.95,
  2.26,    2.26,    2.26,    2.26,
  1.93,    1.93,    1.93,    1.93,
  1.84,    1.84,    1.84,    1.84,
  1.62,    1.62,    1.62,    1.62,
  1.22,    1.22,    1.22,    1.22,
  1.73,    1.73,    1.73,    1.73,
  1.92,    1.92,    1.92,    1.92,
  0.87,    0.87,    0.87,    0.87,
  1.43,    1.43,    1.43,    1.43,
  1.91,    1.91,    1.91,    1.91,
  1.23,    1.23,    1.23,    1.23,
  2.21,    2.21,    2.21,    2.21,
  2,       2,       2,       2,
  1.89,    1.89,    1.89,    1.89,
  2.26,    2.26,    2.26,    2.26,
  1.66,    1.66,    1.66,    1.66,
  2.3,     2.3,     2.3,     2.3,
  2.17,    2.17,    2.17,    2.17,
  2.16,    2.16,    2.16,    2.16,
  2.22,    2.22,    2.22,    2.22,
  2.78,    2.78,    2.78,    2.78,
  2.88,    2.88,    2.88,    2.88,
  2.83,    2.83,    2.83,    2.83,
  3.52,    3.52,    3.52,    3.52,
  2.66,    2.66,    2.66,    2.66,
  2.9,     2.9,     2.9,     2.9,
  2.56,    2.56,    2.56,    2.56,
  2.46,    2.46,    2.46,    2.46,
  2.59,    2.59,    2.59,    2.59,
  1.91,    1.91,    1.91,    1.91,
  2.57,    2.57,    2.57,    2.57,
  2.12,    2.12,    2.12,    2.12,
  1.02,    1.02,    1.02,    1.02,
  1.24,    1.24,    1.24,    1.24,
  0.89,    0.89,    0.89,    0.89,
  1.36,    1.36,    1.36,    1.36,
  1.33,    1.33,    1.33,    1.33,
  1.11,    1.11,    1.11,    1.11,
  1.15,    1.15,    1.15,    1.15,
  1.19,    1.19,    1.19,    1.19,
  1.36,    1.36,    1.36,    1.36,
  0.83,    0.83,    0.83,    0.83,
  0.62,    0.62,    0.62,    0.62,
  0.4,     0.4,     0.4,     0.4,
  0.4,     0.4,     0.4,     0.4,
  1.03,    1.03,    1.03,    1.03,
  1.89,    1.89,    1.89,    1.89,
  1.5,     1.5,     1.5,     1.5,
  1.8,     1.8,     1.8,     1.8,
  1.47,    1.47,    1.47,    1.47,
  1.73,    1.73,    1.73,    1.73,
  1.51,    1.51,    1.51,    1.51,
  1.35,    1.35,    1.35,    1.35,
  1.96,    1.96,    1.96,    1.96,
  1.13,    1.13,    1.13,    1.13,
  1.37,    1.37,    1.37,    1.37,
  1.43,    1.43,    1.43,    1.43,
  0.59,    0.59,    0.59,    0.59,
  1.27,    1.27,    1.27,    1.27,
  1.41,    1.41,    1.41,    1.41,
  1.65,    1.65,    1.65,    1.65,
  2.52,    2.52,    2.52,    2.52,
  2.49,    2.49,    2.49,    2.49,
  2.52,    2.52,    2.52,    2.52,
  2.35,    2.35,    2.35,    2.35,
  2.54,    2.54,    2.54,    2.54,
  2.96,    2.96,    2.96,    2.96,
  3.26,    3.26,    3.26,    3.26,
  3.55,    3.55,    3.55,    3.55,
  3.79,    3.79,    3.79,    3.79,
  3.94,    3.94,    3.94,    3.94,
  4.46,    4.46,    4.46,    4.46,
  4.27,    4.27,    4.27,    4.27,
  4.39,    4.39,    4.39,    4.39,
  3.9,     3.9,     3.9,     3.9,
  4.99,    4.99,    4.99,    4.99,
  4.52,    4.52,    4.52,    4.52,
  4.33,    4.33,    4.33,    4.33,
  4.2,     4.2,     4.2,     4.2,
  4.77,    4.77,    4.77,    4.77,
  4.96,    4.96,    4.96,    4.96,
  4.7,     4.7,     4.7,     4.7,
  3.59,    3.59,    3.59,    3.59,
  4.34,    4.34,    4.34,    4.34,
  3.99,    3.99,    3.99,    3.99,
  3.57,    3.57,    3.57,    3.57,
  2.99,    2.99,    2.99,    2.99,
  2.79,    2.79,    2.79,    2.79,
  3.03,    3.03,    3.03,    3.03,
  3.45,    3.45,    3.45,    3.45,
  3.68,    3.68,    3.68,    3.68,
  3.78,    3.78,    3.78,    3.78,
  3.83,    3.83,    3.83,    3.83,
  4.03,    4.03,    4.03,    4.03,
  3.67,    3.67,    3.67,    3.67,
  3.43,    3.43,    3.43,    3.43,
  3.2,     3.2,     3.2,     3.2,
  3.23,    3.23,    3.23,    3.23,
  3.36,    3.36,    3.36,    3.36,
  3.25,    3.25,    3.25,    3.25,
  2.8,     2.8,     2.8,     2.8,
  2.91,    2.91,    2.91,    2.91,
  2.9,     2.9,     2.9,     2.9,
  2.49,    2.49,    2.49,    2.49,
  2.91,    2.91,    2.91,    2.91,
  2.96,    2.96,    2.96,    2.96,
  2.93,    2.93,    2.93,    2.93,
  3.52,    3.52,    3.52,    3.52,
  3.36,    3.36,    3.36,    3.36,
  3.15,    3.15,    3.15,    3.15,
  3.31,    3.31,    3.31,    3.31,
  3.31,    3.31,    3.31,    3.31,
  3.1,     3.1,     3.1,     3.1,
  2.89,    2.89,    2.89,    2.89,
  2.53,    2.53,    2.53,    2.53,
  3.16,    3.16,    3.16,    3.16,
  3.18,    3.18,    3.18,    3.18,
  3.86,    3.86,    3.86,    3.86,
  3.55,    3.55,    3.55,    3.55,
  3.71,    3.71,    3.71,    3.71,
  4.04,    4.04,    4.04,    4.04,
  3.72,    3.72,    3.72,    3.72,
  3.76,    3.76,    3.76,    3.76,
  3.58,    3.58,    3.58,    3.58,
  2.8,     2.8,     2.8,     2.8,
  2.42,    2.42,    2.42,    2.42,
  2.68,    2.68,    2.68,    2.68,
  2.9,     2.9,     2.9,     2.9,
  3.22,    3.22,    3.22,    3.22,
  2.65,    2.65,    2.65,    2.65,
  2.58,    2.58,    2.58,    2.58,
  2.96,    2.96,    2.96,    2.96,
  2.49,    2.49,    2.49,    2.49,
  2.14,    2.14,    2.14,    2.14,
  2.03,    2.03,    2.03,    2.03,
  1.91,    1.91,    1.91,    1.91,
  2.36,    2.36,    2.36,    2.36,
  2.03,    2.03,    2.03,    2.03,
  1.39,    1.39,    1.39,    1.39,
  0.7,     0.7,     0.7,     0.7,
  1.57,    1.57,    1.57,    1.57,
  1.19,    1.19,    1.19,    1.19,
  0.64,    0.64,    0.64,    0.64,
  0.66,    0.66,    0.66,    0.66,
  0.44,    0.44,    0.44,    0.44,
  1.79,    1.79,    1.79,    1.79,
  1.89,    1.89,    1.89,    1.89,
  1.74,    1.74,    1.74,    1.74,
  2.2,     2.2,     2.2,     2.2,
  0.85,    0.85,    0.85,    0.85,
  1.73,    1.73,    1.73,    1.73,
  1.42,    1.42,    1.42,    1.42,
  1.03,    1.03,    1.03,    1.03,
  1.08,    1.08,    1.08,    1.08,
  0.58,    0.58,    0.58,    0.58,
  0.78,    0.78,    0.78,    0.78,
  1.42,    1.42,    1.42,    1.42,
  2.35,    2.35,    2.35,    2.35,
  1.64,    1.64,    1.64,    1.64,
  2.09,    2.09,    2.09,    2.09,
  2.31,    2.31,    2.31,    2.31,
  2.93,    2.93,    2.93,    2.93,
  2.46,    2.46,    2.46,    2.46,
  2.53,    2.53,    2.53,    2.53,
  2.45,    2.45,    2.45,    2.45,
  2.5,     2.5,     2.5,     2.5,
  2.13,    2.13,    2.13,    2.13,
  2.56,    2.56,    2.56,    2.56,
  2.01,    2.01,    2.01,    2.01,
  1.63,    1.63,    1.63,    1.63,
  2.41,    2.41,    2.41,    2.41,
  2.64,    2.64,    2.64,    2.64,
  2,       2,       2,       2,
  2.18,    2.18,    2.18,    2.18,
  2.06,    2.06,    2.06,    2.06,
  1.76,    1.76,    1.76,    1.76,
  1.88,    1.88,    1.88,    1.88,
  1.25,    1.25,    1.25,    1.25,
  1.23,    1.23,    1.23,    1.23,
  0.83,    0.83,    0.83,    0.83,
  2.52,    2.52,    2.52,    2.52,
  1.22,    1.22,    1.22,    1.22,
  0.82,    0.82,    0.82,    0.82,
  0.23,    0.23,    0.23,    0.23,
  1.01,    1.01,    1.01,    1.01,
  2.09,    2.09,    2.09,    2.09,
  1.95,    1.95,    1.95,    1.95,
  1.88,    1.88,    1.88,    1.88,
  2.57,    2.57,    2.57,    2.57,
  2.35,    2.35,    2.35,    2.35,
  2.53,    2.53,    2.53,    2.53,
  2.32,    2.32,    2.32,    2.32,
  1.78,    1.78,    1.78,    1.78,
  1.76,    1.76,    1.76,    1.76,
  2.2,     2.2,     2.2,     2.2,
  3.12,    3.12,    3.12,    3.12,
  2.54,    2.54,    2.54,    2.54,
  2.62,    2.62,    2.62,    2.62,
  1.79,    1.79,    1.79,    1.79,
  2.03,    2.03,    2.03,    2.03,
  2.02,    2.02,    2.02,    2.02,
  1.4,     1.4,     1.4,     1.4,
  2.6,     2.6,     2.6,     2.6,
  2.35,    2.35,    2.35,    2.35,
  1.85,    1.85,    1.85,    1.85,
  1.71,    1.71,    1.71,    1.71,
  1.4,     1.4,     1.4,     1.4,
  1.65,    1.65,    1.65,    1.65,
  1.79,    1.79,    1.79,    1.79,
  2.85,    2.85,    2.85,    2.85,
  3.57,    3.57,    3.57,    3.57,
  4.06,    4.06,    4.06,    4.06,
  3.83,    3.83,    3.83,    3.83,
  3.9,     3.9,     3.9,     3.9,
  3.58,    3.58,    3.58,    3.58,
  3.43,    3.43,    3.43,    3.43,
  3.7,     3.7,     3.7,     3.7,
  3.26,    3.26,    3.26,    3.26,
  2.73,    2.73,    2.73,    2.73,
  2.66,    2.66,    2.66,    2.66,
  1.98,    1.98,    1.98,    1.98,
  1.8,     1.8,     1.8,     1.8,
  1.56,    1.56,    1.56,    1.56,
  1.23,    1.23,    1.23,    1.23,
  0.64,    0.64,    0.64,    0.64,
  0.4,     0.4,     0.4,     0.4,
  0.53,    0.53,    0.53,    0.53,
  0.26,    0.26,    0.26,    0.26,
  0.19,    0.19,    0.19,    0.19,
  0.68,    0.68,    0.68,    0.68,
  1.09,    1.09,    1.09,    1.09,
  1.36,    1.36,    1.36,    1.36,
  1.28,    1.28,    1.28,    1.28,
  1.13,    1.13,    1.13,    1.13,
  0.82,    0.82,    0.82,    0.82,
  0.33,    0.33,    0.33,    0.33,
  0.52,    0.52,    0.52,    0.52,
  1.1,     1.1,     1.1,     1.1,
  1.27,    1.27,    1.27,    1.27,
  1.4,     1.4,     1.4,     1.4,
  1.69,    1.69,    1.69,    1.69,
  1.63,    1.63,    1.63,    1.63,
  1.89,    1.89,    1.89,    1.89,
  2.12,    2.12,    2.12,    2.12,
  2,       2,       2,       2,
  1.53,    1.53,    1.53,    1.53,
  2.35,    2.35,    2.35,    2.35,
  2.205,   2.205,   2.205,   2.205,
  2.297,   2.297,   2.297,   2.297,
  2.2,     2.2,     2.2,     2.2,
  2.307,   2.307,   2.307,   2.307,
  2.496,   2.496,   2.496,   2.496,
  2.608,   2.608,   2.608,   2.608,
  2.905,   2.905,   2.905,   2.905,
  3.07,    3.07,    3.07,    3.07,
  3.165,   3.165,   3.165,   3.165,
  3.254,   3.254,   3.254,   3.254,
  3.441,   3.441,   3.441,   3.441,
  3.5,     3.5,     3.5,     3.5,
  3.819,   3.819,   3.819,   3.819,
  3.461,   3.461,   3.461,   3.461,
  3.5,     3.5,     3.5,     3.5,
  3.691,   3.691,   3.691,   3.691,
  3.882,   3.882,   3.882,   3.882,
  3.811,   3.811,   3.811,   3.811,
  3.722,   3.722,   3.722,   3.722,
  3.775,   3.775,   3.775,   3.775,
  3.585,   3.585,   3.585,   3.585,
  3.421,   3.421,   3.421,   3.421,
  2.938,   2.938,   2.938,   2.938,
  2.962,   2.962,   2.962,   2.962,
  3.072,   3.072,   3.072,   3.072,
  2.988,   2.988,   2.988,   2.988,
  2.721,   2.721,   2.721,   2.721,
  2.628,   2.628,   2.628,   2.628,
  2.294,   2.294,   2.294,   2.294,
  2.208,   2.208,   2.208,   2.208,
  1.999,   1.999,   1.999,   1.999,
  2.076,   2.076,   2.076,   2.076,
  2.128,   2.128,   2.128,   2.128,
  2.357,   2.357,   2.357,   2.357,
  2.346,   2.346,   2.346,   2.346,
  2.219,   2.219,   2.219,   2.219,
  2.047,   2.047,   2.047,   2.047,
  2.29,    2.29,    2.29,    2.29,
  2.386,   2.386,   2.386,   2.386,
  2.308,   2.308,   2.308,   2.308,
  2.237,   2.237,   2.237,   2.237,
  2.298,   2.298,   2.298,   2.298,
  2.353,   2.353,   2.353,   2.353,
  2.414,   2.414,   2.414,   2.414,
  2.468,   2.468,   2.468,   2.468,
  2.222,   2.222,   2.222,   2.222,
  2.291,   2.291,   2.291,   2.291,
  2.35,    2.35,    2.35,    2.35,
  2.205,   2.205,   2.205,   2.205,
  2.297,   2.297,   2.297,   2.297,
  2.2,     2.2,     2.2,     2.2,
  2.307,   2.307,   2.307,   2.307,
  2.496,   2.496,   2.496,   2.496,
  2.608,   2.608,   2.608,   2.608,
  2.905,   2.905,   2.905,   2.905,
  3.07,    3.07,    3.07,    3.07,
  3.165,   3.165,   3.165,   3.165,
  3.254,   3.254,   3.254,   3.254,
  3.441,   3.441,   3.441,   3.441,
  3.5,     3.5,     3.5,     3.5,
  3.819,   3.819,   3.819,   3.819,
  3.461,   3.461,   3.461,   3.461,
  3.5,     3.5,     3.5,     3.5,
  3.691,   3.691,   3.691,   3.691,
  3.882,   3.882,   3.882,   3.882,
  3.811,   3.811,   3.811,   3.811,
  3.722,   3.722,   3.722,   3.722,
  3.775,   3.775,   3.775,   3.775,
  3.585,   3.585,   3.585,   3.585,
  3.421,   3.421,   3.421,   3.421,
  2.938,   2.938,   2.938,   2.938,
  2.962,   2.962,   2.962,   2.962,
  3.072,   3.072,   3.072,   3.072,
  2.988,   2.988,   2.988,   2.988,
  2.721,   2.721,   2.721,   2.721,
  2.628,   2.628,   2.628,   2.628,
  2.294,   2.294,   2.294,   2.294,
  2.208,   2.208,   2.208,   2.208,
  1.999,   1.999,   1.999,   1.999,
  2.076,   2.076,   2.076,   2.076,
  2.128,   2.128,   2.128,   2.128,
  2.357,   2.357,   2.357,   2.357,
  2.346,   2.346,   2.346,   2.346,
  2.219,   2.219,   2.219,   2.219,
  2.047,   2.047,   2.047,   2.047,
  2.29,    2.29,    2.29,    2.29,
  2.386,   2.386,   2.386,   2.386,
  2.715,   2.715,   2.715,   2.715,
  2.514,   2.514,   2.514,   2.514,
  2.289,   2.289,   2.289,   2.289,
  2.494,   2.494,   2.494,   2.494,
  2.333,   2.333,   2.333,   2.333,
  2.428,   2.428,   2.428,   2.428,
  2.222,   2.222,   2.222,   2.222,
  2.378,   2.378,   2.378,   2.378,
  2.375,   2.375,   2.375,   2.375,
  2.252,   2.252,   2.252,   2.252,
  2.444,   2.444,   2.444,   2.444,
  2.393,   2.393,   2.393,   2.393,
  2.391,   2.391,   2.391,   2.391,
  2.408,   2.408,   2.408,   2.408,
  2.473,   2.473,   2.473,   2.473,
  2.745,   2.745,   2.745,   2.745,
  2.967,   2.967,   2.967,   2.967,
  3.075,   3.075,   3.075,   3.075,
  3.088,   3.088,   3.088,   3.088,
  3.108,   3.108,   3.108,   3.108,
  3.262,   3.262,   3.262,   3.262,
  3.173,   3.173,   3.173,   3.173,
  3.415,   3.415,   3.415,   3.415,
  3.33,    3.33,    3.33,    3.33,
  3.472,   3.472,   3.472,   3.472,
  3.407,   3.407,   3.407,   3.407,
  3.713,   3.713,   3.713,   3.713,
  3.772,   3.772,   3.772,   3.772,
  3.588,   3.588,   3.588,   3.588,
  3.571,   3.571,   3.571,   3.571,
  3.748,   3.748,   3.748,   3.748,
  3.507,   3.507,   3.507,   3.507,
  3.458,   3.458,   3.458,   3.458,
  3.538,   3.538,   3.538,   3.538,
  3.572,   3.572,   3.572,   3.572,
  3.741,   3.741,   3.741,   3.741,
  3.395,   3.395,   3.395,   3.395,
  3.085,   3.085,   3.085,   3.085,
  3.178,   3.178,   3.178,   3.178,
  3.147,   3.147,   3.147,   3.147,
  2.812,   2.812,   2.812,   2.812,
  2.702,   2.702,   2.702,   2.702,
  2.621,   2.621,   2.621,   2.621,
  2.548,   2.548,   2.548,   2.548,
  2.719,   2.719,   2.719,   2.719,
  2.646,   2.646,   2.646,   2.646,
  2.725,   2.725,   2.725,   2.725,
  2.571,   2.571,   2.571,   2.571,
  2.715,   2.715,   2.715,   2.715,
  2.514,   2.514,   2.514,   2.514,
  2.289,   2.289,   2.289,   2.289,
  2.494,   2.494,   2.494,   2.494,
  2.333,   2.333,   2.333,   2.333,
  2.428,   2.428,   2.428,   2.428,
  2.222,   2.222,   2.222,   2.222,
  2.378,   2.378,   2.378,   2.378,
  2.375,   2.375,   2.375,   2.375,
  2.252,   2.252,   2.252,   2.252,
  2.444,   2.444,   2.444,   2.444,
  2.393,   2.393,   2.393,   2.393,
  2.391,   2.391,   2.391,   2.391,
  2.408,   2.408,   2.408,   2.408,
  2.473,   2.473,   2.473,   2.473,
  2.745,   2.745,   2.745,   2.745,
  2.967,   2.967,   2.967,   2.967,
  3.075,   3.075,   3.075,   3.075,
  3.088,   3.088,   3.088,   3.088,
  3.108,   3.108,   3.108,   3.108,
  3.262,   3.262,   3.262,   3.262,
  3.173,   3.173,   3.173,   3.173,
  3.415,   3.415,   3.415,   3.415,
  3.33,    3.33,    3.33,    3.33,
  3.472,   3.472,   3.472,   3.472,
  3.407,   3.407,   3.407,   3.407,
  3.713,   3.713,   3.713,   3.713,
  3.772,   3.772,   3.772,   3.772,
  3.588,   3.588,   3.588,   3.588,
  3.571,   3.571,   3.571,   3.571,
  3.748,   3.748,   3.748,   3.748,
  3.507,   3.507,   3.507,   3.507,
  2.68,    2.68,    2.68,    2.68,
  2.07,    2.07,    2.07,    2.07,
  2.26,    2.26,    2.26,    2.26,
  2.54,    2.54,    2.54,    2.54,
  1.81,    1.81,    1.81,    1.81,
  1.79,    1.79,    1.79,    1.79,
  1.89,    1.89,    1.89,    1.89,
  1.29,    1.29,    1.29,    1.29,
  1.79,    1.79,    1.79,    1.79,
  2.24,    2.24,    2.24,    2.24,
  1.53,    1.53,    1.53,    1.53,
  1.27,    1.27,    1.27,    1.27,
  1.88,    1.88,    1.88,    1.88,
  1.8,     1.8,     1.8,     1.8,
  1.54,    1.54,    1.54,    1.54,
  1.41,    1.41,    1.41,    1.41,
  1.68,    1.68,    1.68,    1.68,
  1.24,    1.24,    1.24,    1.24,
  0.92,    0.92,    0.92,    0.92,
  1.77,    1.77,    1.77,    1.77,
  1.72,    1.72,    1.72,    1.72,
  1.21,    1.21,    1.21,    1.21,
  1.24,    1.24,    1.24,    1.24,
  1.06,    1.06,    1.06,    1.06,
  1.56,    1.56,    1.56,    1.56,
  1.82,    1.82,    1.82,    1.82,
  2.02,    2.02,    2.02,    2.02,
  1.68,    1.68,    1.68,    1.68,
  1.74,    1.74,    1.74,    1.74,
  2.32,    2.32,    2.32,    2.32,
  1.91,    1.91,    1.91,    1.91,
  2.35,    2.35,    2.35,    2.35,
  2.1,     2.1,     2.1,     2.1,
  2.14,    2.14,    2.14,    2.14,
  1.36,    1.36,    1.36,    1.36,
  2.12,    2.12,    2.12,    2.12,
  2.17,    2.17,    2.17,    2.17,
  1.35,    1.35,    1.35,    1.35,
  2.46,    2.46,    2.46,    2.46,
  2.75,    2.75,    2.75,    2.75,
  3.17,    3.17,    3.17,    3.17,
  2.75,    2.75,    2.75,    2.75,
  1.95,    1.95,    1.95,    1.95,
  3.03,    3.03,    3.03,    3.03,
  2.52,    2.52,    2.52,    2.52,
  2.56,    2.56,    2.56,    2.56,
  2.84,    2.84,    2.84,    2.84,
  2.95,    2.95,    2.95,    2.95,
  2.94,    2.94,    2.94,    2.94,
  2.96,    2.96,    2.96,    2.96,
  3.06,    3.06,    3.06,    3.06,
  3.77,    3.77,    3.77,    3.77,
  3.35,    3.35,    3.35,    3.35,
  3.06,    3.06,    3.06,    3.06,
  3.29,    3.29,    3.29,    3.29,
  2.81,    2.81,    2.81,    2.81,
  1.95,    1.95,    1.95,    1.95,
  1.99,    1.99,    1.99,    1.99,
  2.33,    2.33,    2.33,    2.33,
  2.61,    2.61,    2.61,    2.61,
  2.7,     2.7,     2.7,     2.7,
  2.47,    2.47,    2.47,    2.47,
  2.05,    2.05,    2.05,    2.05,
  2.17,    2.17,    2.17,    2.17,
  2.29,    2.29,    2.29,    2.29,
  2.36,    2.36,    2.36,    2.36,
  2.45,    2.45,    2.45,    2.45,
  2.39,    2.39,    2.39,    2.39,
  2.3,     2.3,     2.3,     2.3,
  2.57,    2.57,    2.57,    2.57,
  2.13,    2.13,    2.13,    2.13,
  2.32,    2.32,    2.32,    2.32,
  2.38,    2.38,    2.38,    2.38,
  2.08,    2.08,    2.08,    2.08,
  2.49,    2.49,    2.49,    2.49,
  2.37,    2.37,    2.37,    2.37,
  2.49,    2.49,    2.49,    2.49,
  2.25,    2.25,    2.25,    2.25,
  2.94,    2.94,    2.94,    2.94,
  2.92,    2.92,    2.92,    2.92,
  3.35,    3.35,    3.35,    3.35,
  3.12,    3.12,    3.12,    3.12,
  3.11,    3.11,    3.11,    3.11,
  2.45,    2.45,    2.45,    2.45,
  3.1,     3.1,     3.1,     3.1,
  2.55,    2.55,    2.55,    2.55,
  2.3,     2.3,     2.3,     2.3,
  2.28,    2.28,    2.28,    2.28,
  2.52,    2.52,    2.52,    2.52,
  2.35,    2.35,    2.35,    2.35,
  2.53,    2.53,    2.53,    2.53,
  2.94,    2.94,    2.94,    2.94,
  2.92,    2.92,    2.92,    2.92,
  2.35,    2.35,    2.35,    2.35,
  3.16,    3.16,    3.16,    3.16,
  2.41,    2.41,    2.41,    2.41,
  2.51,    2.51,    2.51,    2.51,
  2.66,    2.66,    2.66,    2.66,
  3.02,    3.02,    3.02,    3.02,
  3.44,    3.44,    3.44,    3.44,
  2.72,    2.72,    2.72,    2.72,
  2.56,    2.56,    2.56,    2.56,
  2.29,    2.29,    2.29,    2.29,
  1.99,    1.99,    1.99,    1.99,
  1.89,    1.89,    1.89,    1.89,
  2.17,    2.17,    2.17,    2.17,
  2.43,    2.43,    2.43,    2.43,
  2.57,    2.57,    2.57,    2.57,
  2.6,     2.6,     2.6,     2.6,
  2.17,    2.17,    2.17,    2.17,
  2.44,    2.44,    2.44,    2.44,
  2.41,    2.41,    2.41,    2.41,
  2.52,    2.52,    2.52,    2.52,
  3.16,    3.16,    3.16,    3.16,
  3.18,    3.18,    3.18,    3.18,
  3.06,    3.06,    3.06,    3.06,
  2.8,     2.8,     2.8,     2.8,
  2.95,    2.95,    2.95,    2.95,
  2.88,    2.88,    2.88,    2.88,
  2.92,    2.92,    2.92,    2.92,
  2.48,    2.48,    2.48,    2.48,
  2.28,    2.28,    2.28,    2.28,
  2.46,    2.46,    2.46,    2.46,
  2.68,    2.68,    2.68,    2.68,
  2.15,    2.15,    2.15,    2.15,
  1.98,    1.98,    1.98,    1.98,
  1.36,    1.36,    1.36,    1.36,
  1.74,    1.74,    1.74,    1.74,
  2.17,    2.17,    2.17,    2.17,
  2.13,    2.13,    2.13,    2.13,
  1.63,    1.63,    1.63,    1.63,
  3.13,    3.13,    3.13,    3.13,
  3.07,    3.07,    3.07,    3.07,
  2.81,    2.81,    2.81,    2.81,
  2.94,    2.94,    2.94,    2.94,
  1.72,    1.72,    1.72,    1.72,
  1.56,    1.56,    1.56,    1.56,
  1.86,    1.86,    1.86,    1.86,
  2.08,    2.08,    2.08,    2.08,
  2.69,    2.69,    2.69,    2.69,
  2.14,    2.14,    2.14,    2.14,
  2.21,    2.21,    2.21,    2.21,
  2.06,    2.06,    2.06,    2.06,
  2.47,    2.47,    2.47,    2.47,
  2.16,    2.16,    2.16,    2.16,
  2.62,    2.62,    2.62,    2.62,
  2.63,    2.63,    2.63,    2.63,
  2.78,    2.78,    2.78,    2.78,
  2.27,    2.27,    2.27,    2.27,
  2.58,    2.58,    2.58,    2.58,
  2.89,    2.89,    2.89,    2.89,
  3.99,    3.99,    3.99,    3.99,
  3.52,    3.52,    3.52,    3.52,
  2.88,    2.88,    2.88,    2.88,
  3.22,    3.22,    3.22,    3.22,
  3,       3,       3,       3,
  2.78,    2.78,    2.78,    2.78,
  2.74,    2.74,    2.74,    2.74,
  2.78,    2.78,    2.78,    2.78,
  2.41,    2.41,    2.41,    2.41,
  2.33,    2.33,    2.33,    2.33,
  1.98,    1.98,    1.98,    1.98,
  1.59,    1.59,    1.59,    1.59,
  1.97,    1.97,    1.97,    1.97,
  1.85,    1.85,    1.85,    1.85,
  1.68,    1.68,    1.68,    1.68,
  1.2,     1.2,     1.2,     1.2,
  1.66,    1.66,    1.66,    1.66,
  1.87,    1.87,    1.87,    1.87,
  0.67,    0.67,    0.67,    0.67,
  1.03,    1.03,    1.03,    1.03,
  1.15,    1.15,    1.15,    1.15,
  1.34,    1.34,    1.34,    1.34,
  1,       1,       1,       1,
  1.42,    1.42,    1.42,    1.42,
  1.54,    1.54,    1.54,    1.54,
  0.75,    0.75,    0.75,    0.75,
  1.4,     1.4,     1.4,     1.4,
  0.95,    0.95,    0.95,    0.95,
  0.77,    0.77,    0.77,    0.77,
  1.23,    1.23,    1.23,    1.23,
  1.52,    1.52,    1.52,    1.52,
  1.92,    1.92,    1.92,    1.92,
  2.06,    2.06,    2.06,    2.06,
  1.54,    1.54,    1.54,    1.54,
  1.6,     1.6,     1.6,     1.6,
  3.713,   3.713,   3.713,   3.713,
  2.59,    2.59,    2.59,    2.59,
  2.53,    2.53,    2.53,    2.53,
  3.07,    3.07,    3.07,    3.07,
  2.98,    2.98,    2.98,    2.98,
  3.89,    3.89,    3.89,    3.89,
  3.32,    3.32,    3.32,    3.32,
  3.95,    3.95,    3.95,    3.95,
  4.01,    4.01,    4.01,    4.01,
  4.14,    4.14,    4.14,    4.14,
  3.68,    3.68,    3.68,    3.68,
  2.87,    2.87,    2.87,    2.87,
  3.22,    3.22,    3.22,    3.22,
  3.46,    3.46,    3.46,    3.46,
  3.46,    3.46,    3.46,    3.46,
  3.77,    3.77,    3.77,    3.77,
  3.4,     3.4,     3.4,     3.4,
  3.7,     3.7,     3.7,     3.7,
  3.76,    3.76,    3.76,    3.76,
  2.87,    2.87,    2.87,    2.87,
  2.95,    2.95,    2.95,    2.95,
  2.78,    2.78,    2.78,    2.78,
  2.72,    2.72,    2.72,    2.72,
  2.54,    2.54,    2.54,    2.54,
  1.84,    1.84,    1.84,    1.84,
  2.25,    2.25,    2.25,    2.25,
  2.25,    2.25,    2.25,    2.25,
  2.9,     2.9,     2.9,     2.9,
  2.78,    2.78,    2.78,    2.78,
  3.14,    3.14,    3.14,    3.14,
  2.84,    2.84,    2.84,    2.84,
  2.82,    2.82,    2.82,    2.82,
  3.12,    3.12,    3.12,    3.12,
  2.75,    2.75,    2.75,    2.75,
  3.25,    3.25,    3.25,    3.25,
  2.31,    2.31,    2.31,    2.31,
  2.17,    2.17,    2.17,    2.17,
  2.55,    2.55,    2.55,    2.55,
  2.63,    2.63,    2.63,    2.63,
  2.49,    2.49,    2.49,    2.49,
  2.88,    2.88,    2.88,    2.88,
  3.24,    3.24,    3.24,    3.24,
  3.59,    3.59,    3.59,    3.59,
  2.66,    2.66,    2.66,    2.66,
  2.88,    2.88,    2.88,    2.88,
  3.02,    3.02,    3.02,    3.02,
  3.38,    3.38,    3.38,    3.38,
  3.41,    3.41,    3.41,    3.41,
  3.37,    3.37,    3.37,    3.37,
  3.66,    3.66,    3.66,    3.66,
  3.85,    3.85,    3.85,    3.85,
  3.36,    3.36,    3.36,    3.36,
  4.65,    4.65,    4.65,    4.65,
  3.99,    3.99,    3.99,    3.99,
  3.31,    3.31,    3.31,    3.31,
  3.77,    3.77,    3.77,    3.77,
  4.15,    4.15,    4.15,    4.15,
  4.21,    4.21,    4.21,    4.21,
  3.87,    3.87,    3.87,    3.87,
  3.56,    3.56,    3.56,    3.56,
  3.51,    3.51,    3.51,    3.51,
  3.9,     3.9,     3.9,     3.9,
  3.05,    3.05,    3.05,    3.05,
  2.26,    2.26,    2.26,    2.26,
  2.25,    2.25,    2.25,    2.25,
  2.18,    2.18,    2.18,    2.18,
  1.85,    1.85,    1.85,    1.85,
  1.95,    1.95,    1.95,    1.95,
  2.31,    2.31,    2.31,    2.31,
  1.86,    1.86,    1.86,    1.86,
  2.89,    2.89,    2.89,    2.89,
  2.85,    2.85,    2.85,    2.85,
  1.96,    1.96,    1.96,    1.96,
  2.12,    2.12,    2.12,    2.12,
  2.12,    2.12,    2.12,    2.12,
  1.83,    1.83,    1.83,    1.83,
  1.45,    1.45,    1.45,    1.45,
  2.45,    2.45,    2.45,    2.45,
  2.28,    2.28,    2.28,    2.28,
  1.72,    1.72,    1.72,    1.72,
  1.78,    1.78,    1.78,    1.78,
  2.04,    2.04,    2.04,    2.04,
  2.11,    2.11,    2.11,    2.11,
  2.65,    2.65,    2.65,    2.65,
  2.91,    2.91,    2.91,    2.91,
  3.04,    3.04,    3.04,    3.04,
  2.89,    2.89,    2.89,    2.89,
  2.82,    2.82,    2.82,    2.82,
  3.12,    3.12,    3.12,    3.12,
  2.85,    2.85,    2.85,    2.85,
  2.54,    2.54,    2.54,    2.54,
  1.95,    1.95,    1.95,    1.95,
  2.37,    2.37,    2.37,    2.37,
  1.93,    1.93,    1.93,    1.93,
  2.37,    2.37,    2.37,    2.37,
  2.28,    2.28,    2.28,    2.28,
  2.44,    2.44,    2.44,    2.44,
  2.2,     2.2,     2.2,     2.2,
  2.31,    2.31,    2.31,    2.31,
  2.34,    2.34,    2.34,    2.34,
  2.94,    2.94,    2.94,    2.94,
  3.29,    3.29,    3.29,    3.29,
  3.64,    3.64,    3.64,    3.64,
  2.34,    2.34,    2.34,    2.34,
  2.21,    2.21,    2.21,    2.21,
  2.6,     2.6,     2.6,     2.6,
  2.17,    2.17,    2.17,    2.17,
  2.71,    2.71,    2.71,    2.71,
  2.56,    2.56,    2.56,    2.56,
  3.03,    3.03,    3.03,    3.03,
  2.36,    2.36,    2.36,    2.36,
  2.06,    2.06,    2.06,    2.06,
  2.13,    2.13,    2.13,    2.13,
  1.98,    1.98,    1.98,    1.98,
  2.13,    2.13,    2.13,    2.13,
  2.22,    2.22,    2.22,    2.22,
  2.2,     2.2,     2.2,     2.2,
  1.87,    1.87,    1.87,    1.87,
  2.1,     2.1,     2.1,     2.1,
  2.1,     2.1,     2.1,     2.1,
  1.87,    1.87,    1.87,    1.87,
  1.84,    1.84,    1.84,    1.84,
  1.63,    1.63,    1.63,    1.63,
  1.41,    1.41,    1.41,    1.41,
  1.67,    1.67,    1.67,    1.67,
  1.57,    1.57,    1.57,    1.57,
  1.83,    1.83,    1.83,    1.83,
  1.58,    1.58,    1.58,    1.58,
  2.11,    2.11,    2.11,    2.11,
  1.42,    1.42,    1.42,    1.42,
  1.24,    1.24,    1.24,    1.24,
  1.26,    1.26,    1.26,    1.26,
  0.63,    0.63,    0.63,    0.63,
  0.83,    0.83,    0.83,    0.83,
  1.39,    1.39,    1.39,    1.39,
  1.44,    1.44,    1.44,    1.44,
  1.85,    1.85,    1.85,    1.85,
  1.12,    1.12,    1.12,    1.12,
  1.62,    1.62,    1.62,    1.62,
  1.4,     1.4,     1.4,     1.4,
  1.78,    1.78,    1.78,    1.78,
  2.42,    2.42,    2.42,    2.42,
  2.76,    2.76,    2.76,    2.76,
  3.31,    3.31,    3.31,    3.31,
  2.38,    2.38,    2.38,    2.38,
  3.18,    3.18,    3.18,    3.18,
  2.94,    2.94,    2.94,    2.94,
  2.92,    2.92,    2.92,    2.92,
  3.23,    3.23,    3.23,    3.23,
  2.41,    2.41,    2.41,    2.41,
  3.13,    3.13,    3.13,    3.13,
  3.67,    3.67,    3.67,    3.67,
  3.72,    3.72,    3.72,    3.72,
  3.92,    3.92,    3.92,    3.92,
  3.02,    3.02,    3.02,    3.02,
  2.36,    2.36,    2.36,    2.36,
  2.9,     2.9,     2.9,     2.9,
  2.96,    2.96,    2.96,    2.96,
  2.69,    2.69,    2.69,    2.69,
  2.12,    2.12,    2.12,    2.12,
  1.83,    1.83,    1.83,    1.83,
  2.08,    2.08,    2.08,    2.08,
  2.05,    2.05,    2.05,    2.05,
  2.19,    2.19,    2.19,    2.19,
  2.23,    2.23,    2.23,    2.23,
  2.17,    2.17,    2.17,    2.17,
  2.715,   2.715,   2.715,   2.715,
  1.63,    1.63,    1.63,    1.63,
  2.11,    2.11,    2.11,    2.11,
  2.15,    2.15,    2.15,    2.15,
  0.85,    0.85,    0.85,    0.85,
  1.14,    1.14,    1.14,    1.14,
  0.57,    0.57,    0.57,    0.57,
  1.28,    1.28,    1.28,    1.28,
  1.72,    1.72,    1.72,    1.72,
  1.95,    1.95,    1.95,    1.95,
  2.3,     2.3,     2.3,     2.3,
  2.45,    2.45,    2.45,    2.45,
  2.18,    2.18,    2.18,    2.18,
  2.49,    2.49,    2.49,    2.49,
  2.79,    2.79,    2.79,    2.79,
  2.44,    2.44,    2.44,    2.44,
  2.69,    2.69,    2.69,    2.69,
  2.96,    2.96,    2.96,    2.96,
  3,       3,       3,       3,
  2.42,    2.42,    2.42,    2.42,
  2.69,    2.69,    2.69,    2.69,
  3.24,    3.24,    3.24,    3.24,
  3.1,     3.1,     3.1,     3.1,
  3.28,    3.28,    3.28,    3.28,
  3.01,    3.01,    3.01,    3.01,
  2.54,    2.54,    2.54,    2.54,
  3.89,    3.89,    3.89,    3.89,
  3.67,    3.67,    3.67,    3.67,
  3.29,    3.29,    3.29,    3.29,
  2.66,    2.66,    2.66,    2.66,
  2.87,    2.87,    2.87,    2.87,
  2.81,    2.81,    2.81,    2.81,
  2.01,    2.01,    2.01,    2.01,
  2.77,    2.77,    2.77,    2.77,
  2.85,    2.85,    2.85,    2.85,
  2.95,    2.95,    2.95,    2.95,
  3.33,    3.33,    3.33,    3.33,
  3.36,    3.36,    3.36,    3.36,
  3.08,    3.08,    3.08,    3.08,
  3.1,     3.1,     3.1,     3.1,
  2.34,    2.34,    2.34,    2.34,
  2.35,    2.35,    2.35,    2.35,
  2.54,    2.54,    2.54,    2.54,
  2.63,    2.63,    2.63,    2.63,
  2.26,    2.26,    2.26,    2.26,
  2.61,    2.61,    2.61,    2.61,
  2.7,     2.7,     2.7,     2.7,
  2.9,     2.9,     2.9,     2.9,
  2.96,    2.96,    2.96,    2.96,
  2.52,    2.52,    2.52,    2.52,
  2.52,    2.52,    2.52,    2.52,
  2.8,     2.8,     2.8,     2.8,
  2.75,    2.75,    2.75,    2.75,
  2.77,    2.77,    2.77,    2.77,
  2.92,    2.92,    2.92,    2.92,
  2.89,    2.89,    2.89,    2.89,
  2.58,    2.58,    2.58,    2.58,
  2.69,    2.69,    2.69,    2.69,
  2.63,    2.63,    2.63,    2.63,
  2.63,    2.63,    2.63,    2.63,
  2.86,    2.86,    2.86,    2.86,
  2.89,    2.89,    2.89,    2.89,
  2.49,    2.49,    2.49,    2.49,
  3.35,    3.35,    3.35,    3.35,
  3.53,    3.53,    3.53,    3.53,
  3.46,    3.46,    3.46,    3.46,
  4.3,     4.3,     4.3,     4.3,
  4.08,    4.08,    4.08,    4.08,
  3.52,    3.52,    3.52,    3.52,
  3.87,    3.87,    3.87,    3.87,
  4.64,    4.64,    4.64,    4.64,
  4.36,    4.36,    4.36,    4.36,
  4.43,    4.43,    4.43,    4.43,
  4,       4,       4,       4,
  4.33,    4.33,    4.33,    4.33,
  5.09,    5.09,    5.09,    5.09,
  4.4,     4.4,     4.4,     4.4,
  4.97,    4.97,    4.97,    4.97,
  5.17,    5.17,    5.17,    5.17,
  4.24,    4.24,    4.24,    4.24,
  4.94,    4.94,    4.94,    4.94,
  4.79,    4.79,    4.79,    4.79,
  4.82,    4.82,    4.82,    4.82,
  5.1,     5.1,     5.1,     5.1,
  4.74,    4.74,    4.74,    4.74,
  4.26,    4.26,    4.26,    4.26,
  3.7,     3.7,     3.7,     3.7,
  3.6,     3.6,     3.6,     3.6,
  3.36,    3.36,    3.36,    3.36,
  2.96,    2.96,    2.96,    2.96,
  2.71,    2.71,    2.71,    2.71,
  2.72,    2.72,    2.72,    2.72,
  3.97,    3.97,    3.97,    3.97,
  3.74,    3.74,    3.74,    3.74,
  3.99,    3.99,    3.99,    3.99,
  3.89,    3.89,    3.89,    3.89,
  3.37,    3.37,    3.37,    3.37,
  3.35,    3.35,    3.35,    3.35,
  2.8,     2.8,     2.8,     2.8,
  3.04,    3.04,    3.04,    3.04,
  3.28,    3.28,    3.28,    3.28,
  2.96,    2.96,    2.96,    2.96,
  2.78,    2.78,    2.78,    2.78,
  2.67,    2.67,    2.67,    2.67,
  2.42,    2.42,    2.42,    2.42,
  2.95,    2.95,    2.95,    2.95,
  3.05,    3.05,    3.05,    3.05,
  2.89,    2.89,    2.89,    2.89,
  3.59,    3.59,    3.59,    3.59,
  3.52,    3.52,    3.52,    3.52,
  4.43,    4.43,    4.43,    4.43,
  4.83,    4.83,    4.83,    4.83,
  5.58,    5.58,    5.58,    5.58,
  5.98,    5.98,    5.98,    5.98,
  6.29,    6.29,    6.29,    6.29,
  6.18,    6.18,    6.18,    6.18,
  5.69,    5.69,    5.69,    5.69,
  6.68,    6.68,    6.68,    6.68,
  6.49,    6.49,    6.49,    6.49,
  6.14,    6.14,    6.14,    6.14,
  6.34,    6.34,    6.34,    6.34,
  6.57,    6.57,    6.57,    6.57,
  7.44,    7.44,    7.44,    7.44,
  6.56,    6.56,    6.56,    6.56,
  6.53,    6.53,    6.53,    6.53,
  7.54,    7.54,    7.54,    7.54,
  7.15,    7.15,    7.15,    7.15,
  6.84,    6.84,    6.84,    6.84,
  6.72,    6.72,    6.72,    6.72,
  7.31,    7.31,    7.31,    7.31,
  6.58,    6.58,    6.58,    6.58,
  6.7,     6.7,     6.7,     6.7,
  6.37,    6.37,    6.37,    6.37,
  5.21,    5.21,    5.21,    5.21,
  6.62,    6.62,    6.62,    6.62,
  5.54,    5.54,    5.54,    5.54,
  5.17,    5.17,    5.17,    5.17,
  5.55,    5.55,    5.55,    5.55,
  3.94,    3.94,    3.94,    3.94,
  3.19,    3.19,    3.19,    3.19,
  4.3,     4.3,     4.3,     4.3,
  4.66,    4.66,    4.66,    4.66,
  4.95,    4.95,    4.95,    4.95,
  4.39,    4.39,    4.39,    4.39,
  4.1,     4.1,     4.1,     4.1,
  3.95,    3.95,    3.95,    3.95,
  3.66,    3.66,    3.66,    3.66,
  3.89,    3.89,    3.89,    3.89,
  4.1,     4.1,     4.1,     4.1,
  4.51,    4.51,    4.51,    4.51,
  4.14,    4.14,    4.14,    4.14,
  3.75,    3.75,    3.75,    3.75,
  3.88,    3.88,    3.88,    3.88,
  3.85,    3.85,    3.85,    3.85,
  3.73,    3.73,    3.73,    3.73,
  4.42,    4.42,    4.42,    4.42,
  3.93,    3.93,    3.93,    3.93,
  4.11,    4.11,    4.11,    4.11,
  4.27,    4.27,    4.27,    4.27,
  4.16,    4.16,    4.16,    4.16,
  5.05,    5.05,    5.05,    5.05,
  4.81,    4.81,    4.81,    4.81,
  5,       5,       5,       5,
  5.4,     5.4,     5.4,     5.4,
  5.56,    5.56,    5.56,    5.56,
  5.37,    5.37,    5.37,    5.37,
  5.82,    5.82,    5.82,    5.82,
  5.9,     5.9,     5.9,     5.9,
  6.49,    6.49,    6.49,    6.49,
  6.38,    6.38,    6.38,    6.38,
  6.22,    6.22,    6.22,    6.22,
  6.37,    6.37,    6.37,    6.37,
  5.36,    5.36,    5.36,    5.36,
  4.86,    4.86,    4.86,    4.86,
  4.97,    4.97,    4.97,    4.97,
  4.31,    4.31,    4.31,    4.31,
  4.62,    4.62,    4.62,    4.62,
  4.69,    4.69,    4.69,    4.69,
  4.47,    4.47,    4.47,    4.47,
  3.93,    3.93,    3.93,    3.93,
  4.6,     4.6,     4.6,     4.6,
  3.47,    3.47,    3.47,    3.47,
  3.47,    3.47,    3.47,    3.47,
  3.41,    3.41,    3.41,    3.41,
  3.18,    3.18,    3.18,    3.18,
  2.83,    2.83,    2.83,    2.83,
  3.03,    3.03,    3.03,    3.03,
  2.5,     2.5,     2.5,     2.5,
  2.63,    2.63,    2.63,    2.63,
  2.54,    2.54,    2.54,    2.54,
  2.91,    2.91,    2.91,    2.91,
  2.94,    2.94,    2.94,    2.94,
  2.91,    2.91,    2.91,    2.91,
  2.49,    2.49,    2.49,    2.49,
  2.57,    2.57,    2.57,    2.57,
  2.65,    2.65,    2.65,    2.65,
  2.35,    2.35,    2.35,    2.35,
  3.2,     3.2,     3.2,     3.2,
  2.9,     2.9,     2.9,     2.9,
  2.83,    2.83,    2.83,    2.83,
  2.66,    2.66,    2.66,    2.66,
  2.61,    2.61,    2.61,    2.61,
  2.61,    2.61,    2.61,    2.61,
  2.24,    2.24,    2.24,    2.24,
  1.81,    1.81,    1.81,    1.81,
  2.12,    2.12,    2.12,    2.12,
  2.36,    2.36,    2.36,    2.36,
  3.19,    3.19,    3.19,    3.19,
  3.47,    3.47,    3.47,    3.47,
  4.15,    4.15,    4.15,    4.15,
  3.57,    3.57,    3.57,    3.57,
  3.53,    3.53,    3.53,    3.53,
  4.36,    4.36,    4.36,    4.36,
  4.68,    4.68,    4.68,    4.68,
  4.28,    4.28,    4.28,    4.28,
  4.1,     4.1,     4.1,     4.1,
  4.09,    4.09,    4.09,    4.09,
  3.83,    3.83,    3.83,    3.83,
  4.21,    4.21,    4.21,    4.21,
  3.28,    3.28,    3.28,    3.28,
  4.27,    4.27,    4.27,    4.27,
  4.01,    4.01,    4.01,    4.01,
  2.96,    2.96,    2.96,    2.96,
  2.48,    2.48,    2.48,    2.48,
  2.97,    2.97,    2.97,    2.97,
  2.39,    2.39,    2.39,    2.39,
  2.66,    2.66,    2.66,    2.66,
  2.55,    2.55,    2.55,    2.55,
  2.21,    2.21,    2.21,    2.21,
  2.31,    2.31,    2.31,    2.31,
  1.9,     1.9,     1.9,     1.9,
  1.83,    1.83,    1.83,    1.83,
  1.79,    1.79,    1.79,    1.79,
  1.95,    1.95,    1.95,    1.95,
  2.73,    2.73,    2.73,    2.73,
  2.7,     2.7,     2.7,     2.7,
  2.44,    2.44,    2.44,    2.44,
  2.44,    2.44,    2.44,    2.44,
  2.38,    2.38,    2.38,    2.38,
  2.22,    2.22,    2.22,    2.22,
  2.62,    2.62,    2.62,    2.62,
  2.79,    2.79,    2.79,    2.79,
  2.86,    2.86,    2.86,    2.86,
  3.06,    3.06,    3.06,    3.06,
  2.48,    2.48,    2.48,    2.48,
  2.15,    2.15,    2.15,    2.15,
  2.55,    2.55,    2.55,    2.55,
  2.51,    2.51,    2.51,    2.51,
  2.57,    2.57,    2.57,    2.57,
  1.09,    1.09,    1.09,    1.09,
  1.71,    1.71,    1.71,    1.71,
  1.18,    1.18,    1.18,    1.18,
  1.2,     1.2,     1.2,     1.2,
  1.25,    1.25,    1.25,    1.25,
  1.18,    1.18,    1.18,    1.18,
  1.22,    1.22,    1.22,    1.22,
  1.24,    1.24,    1.24,    1.24,
  1.56,    1.56,    1.56,    1.56,
  1.15,    1.15,    1.15,    1.15,
  1.06,    1.06,    1.06,    1.06,
  1.01,    1.01,    1.01,    1.01,
  1.45,    1.45,    1.45,    1.45,
  1.38,    1.38,    1.38,    1.38,
  1.22,    1.22,    1.22,    1.22,
  0.92,    0.92,    0.92,    0.92,
  1.18,    1.18,    1.18,    1.18,
  1.06,    1.06,    1.06,    1.06,
  1.38,    1.38,    1.38,    1.38,
  1.94,    1.94,    1.94,    1.94,
  2.35,    2.35,    2.35,    2.35,
  1.22,    1.22,    1.22,    1.22,
  2.11,    2.11,    2.11,    2.11,
  1.96,    1.96,    1.96,    1.96,
  1.41,    1.41,    1.41,    1.41,
  1.49,    1.49,    1.49,    1.49,
  2.02,    2.02,    2.02,    2.02,
  2.99,    2.99,    2.99,    2.99,
  3.07,    3.07,    3.07,    3.07,
  2.81,    2.81,    2.81,    2.81,
  2.03,    2.03,    2.03,    2.03,
  1.76,    1.76,    1.76,    1.76,
  2.19,    2.19,    2.19,    2.19,
  2.29,    2.29,    2.29,    2.29,
  2.45,    2.45,    2.45,    2.45,
  2.65,    2.65,    2.65,    2.65,
  2.66,    2.66,    2.66,    2.66,
  3.23,    3.23,    3.23,    3.23,
  3.21,    3.21,    3.21,    3.21,
  3.3,     3.3,     3.3,     3.3,
  3.16,    3.16,    3.16,    3.16,
  3.15,    3.15,    3.15,    3.15,
  3.43,    3.43,    3.43,    3.43,
  2.69,    2.69,    2.69,    2.69,
  2.92,    2.92,    2.92,    2.92,
  2.82,    2.82,    2.82,    2.82,
  2.92,    2.92,    2.92,    2.92,
  2.71,    2.71,    2.71,    2.71,
  2.98,    2.98,    2.98,    2.98,
  2.96,    2.96,    2.96,    2.96,
  3.44,    3.44,    3.44,    3.44,
  3.08,    3.08,    3.08,    3.08,
  2.37,    2.37,    2.37,    2.37,
  2.25,    2.25,    2.25,    2.25,
  2.16,    2.16,    2.16,    2.16,
  1.59,    1.59,    1.59,    1.59,
  2.12,    2.12,    2.12,    2.12,
  2.45,    2.45,    2.45,    2.45,
  2.98,    2.98,    2.98,    2.98,
  3.67,    3.67,    3.67,    3.67,
  3.87,    3.87,    3.87,    3.87,
  4.08,    4.08,    4.08,    4.08,
  4.18,    4.18,    4.18,    4.18,
  4.21,    4.21,    4.21,    4.21,
  3.95,    3.95,    3.95,    3.95,
  3.93,    3.93,    3.93,    3.93,
  4.22,    4.22,    4.22,    4.22,
  4.65,    4.65,    4.65,    4.65,
  4.95,    4.95,    4.95,    4.95,
  3.95,    3.95,    3.95,    3.95,
  3.86,    3.86,    3.86,    3.86,
  3.96,    3.96,    3.96,    3.96,
  4.36,    4.36,    4.36,    4.36,
  4.59,    4.59,    4.59,    4.59,
  4.27,    4.27,    4.27,    4.27,
  4.25,    4.25,    4.25,    4.25,
  3.85,    3.85,    3.85,    3.85,
  3.72,    3.72,    3.72,    3.72,
  3.29,    3.29,    3.29,    3.29,
  2.79,    2.79,    2.79,    2.79,
  2.69,    2.69,    2.69,    2.69,
  2.67,    2.67,    2.67,    2.67,
  2.88,    2.88,    2.88,    2.88,
  2.97,    2.97,    2.97,    2.97,
  3.06,    3.06,    3.06,    3.06,
  3.11,    3.11,    3.11,    3.11,
  3.08,    3.08,    3.08,    3.08,
  2.85,    2.85,    2.85,    2.85,
  2.98,    2.98,    2.98,    2.98,
  3.08,    3.08,    3.08,    3.08,
  3.07,    3.07,    3.07,    3.07,
  3.17,    3.17,    3.17,    3.17,
  3.01,    3.01,    3.01,    3.01,
  2.67,    2.67,    2.67,    2.67,
  2.81,    2.81,    2.81,    2.81,
  3.08,    3.08,    3.08,    3.08,
  3.29,    3.29,    3.29,    3.29,
  2.89,    2.89,    2.89,    2.89,
  2.68,    2.68,    2.68,    2.68,
  2.4,     2.4,     2.4,     2.4,
  2.12,    2.12,    2.12,    2.12,
  2.43,    2.43,    2.43,    2.43,
  2.16,    2.16,    2.16,    2.16,
  2.53,    2.53,    2.53,    2.53,
  2.7,     2.7,     2.7,     2.7,
  2.52,    2.52,    2.52,    2.52,
  1.99,    1.99,    1.99,    1.99,
  1.58,    1.58,    1.58,    1.58,
  2.12,    2.12,    2.12,    2.12,
  2.72,    2.72,    2.72,    2.72,
  2.82,    2.82,    2.82,    2.82,
  3.83,    3.83,    3.83,    3.83,
  3.54,    3.54,    3.54,    3.54,
  4.62,    4.62,    4.62,    4.62,
  4.64,    4.64,    4.64,    4.64,
  3.8,     3.8,     3.8,     3.8,
  4.28,    4.28,    4.28,    4.28,
  3.69,    3.69,    3.69,    3.69,
  4.04,    4.04,    4.04,    4.04,
  4.13,    4.13,    4.13,    4.13,
  3.37,    3.37,    3.37,    3.37,
  3.59,    3.59,    3.59,    3.59,
  3.42,    3.42,    3.42,    3.42,
  3.41,    3.41,    3.41,    3.41,
  3.29,    3.29,    3.29,    3.29,
  3.35,    3.35,    3.35,    3.35,
  2.13,    2.13,    2.13,    2.13,
  1.94,    1.94,    1.94,    1.94,
  2.08,    2.08,    2.08,    2.08,
  2.22,    2.22,    2.22,    2.22,
  2.17,    2.17,    2.17,    2.17,
  1.9,     1.9,     1.9,     1.9,
  2.29,    2.29,    2.29,    2.29,
  2.41,    2.41,    2.41,    2.41,
  2.37,    2.37,    2.37,    2.37,
  2.75,    2.75,    2.75,    2.75,
  2.71,    2.71,    2.71,    2.71,
  2.76,    2.76,    2.76,    2.76,
  2.6,     2.6,     2.6,     2.6,
  2.44,    2.44,    2.44,    2.44,
  2.61,    2.61,    2.61,    2.61,
  2.79,    2.79,    2.79,    2.79,
  2.93,    2.93,    2.93,    2.93,
  3.11,    3.11,    3.11,    3.11,
  3.11,    3.11,    3.11,    3.11,
  3.13,    3.13,    3.13,    3.13,
  3.5,     3.5,     3.5,     3.5,
  3.65,    3.65,    3.65,    3.65,
  3.7,     3.7,     3.7,     3.7,
  3.61,    3.61,    3.61,    3.61,
  4.29,    4.29,    4.29,    4.29,
  4.41,    4.41,    4.41,    4.41,
  4.49,    4.49,    4.49,    4.49,
  4.67,    4.67,    4.67,    4.67,
  3.95,    3.95,    3.95,    3.95,
  4.35,    4.35,    4.35,    4.35,
  4.76,    4.76,    4.76,    4.76,
  5.2,     5.2,     5.2,     5.2,
  4.19,    4.19,    4.19,    4.19,
  4.35,    4.35,    4.35,    4.35,
  4.61,    4.61,    4.61,    4.61,
  4.28,    4.28,    4.28,    4.28,
  4.51,    4.51,    4.51,    4.51,
  5.22,    5.22,    5.22,    5.22,
  3.71,    3.71,    3.71,    3.71,
  4.52,    4.52,    4.52,    4.52,
  4.35,    4.35,    4.35,    4.35,
  1.23,    1.23,    1.23,    1.23,
  2.74,    2.74,    2.74,    2.74,
  0.63,    0.63,    0.63,    0.63,
  0.77,    0.77,    0.77,    0.77,
  1.29,    1.29,    1.29,    1.29,
  1.19,    1.19,    1.19,    1.19,
  0.87,    0.87,    0.87,    0.87,
  0.58,    0.58,    0.58,    0.58,
  1.15,    1.15,    1.15,    1.15,
  0.59,    0.59,    0.59,    0.59,
  1.21,    1.21,    1.21,    1.21,
  1.81,    1.81,    1.81,    1.81,
  1.49,    1.49,    1.49,    1.49,
  2.26,    2.26,    2.26,    2.26,
  1.73,    1.73,    1.73,    1.73,
  0.77,    0.77,    0.77,    0.77,
  0.86,    0.86,    0.86,    0.86,
  0.26,    0.26,    0.26,    0.26,
  1.33,    1.33,    1.33,    1.33,
  1.26,    1.26,    1.26,    1.26,
  1.59,    1.59,    1.59,    1.59,
  2.15,    2.15,    2.15,    2.15,
  1.9,     1.9,     1.9,     1.9,
  1.52,    1.52,    1.52,    1.52,
  2.13,    2.13,    2.13,    2.13,
  2.14,    2.14,    2.14,    2.14,
  1.88,    1.88,    1.88,    1.88,
  2.38,    2.38,    2.38,    2.38,
  2.03,    2.03,    2.03,    2.03,
  1.54,    1.54,    1.54,    1.54,
  2.35,    2.35,    2.35,    2.35,
  2.26,    2.26,    2.26,    2.26,
  2.1,     2.1,     2.1,     2.1,
  2,       2,       2,       2,
  2.72,    2.72,    2.72,    2.72,
  2.36,    2.36,    2.36,    2.36,
  1.56,    1.56,    1.56,    1.56,
  1.16,    1.16,    1.16,    1.16,
  1.54,    1.54,    1.54,    1.54,
  1.58,    1.58,    1.58,    1.58,
  1.67,    1.67,    1.67,    1.67,
  0.51,    0.51,    0.51,    0.51,
  0.28,    0.28,    0.28,    0.28,
  1.56,    1.56,    1.56,    1.56,
  1.19,    1.19,    1.19,    1.19,
  0.91,    0.91,    0.91,    0.91,
  1.9,     1.9,     1.9,     1.9,
  1.74,    1.74,    1.74,    1.74,
  1.62,    1.62,    1.62,    1.62,
  1.25,    1.25,    1.25,    1.25,
  3.19,    3.19,    3.19,    3.19,
  2.85,    2.85,    2.85,    2.85,
  2.79,    2.79,    2.79,    2.79,
  2.82,    2.82,    2.82,    2.82,
  2.54,    2.54,    2.54,    2.54,
  1.12,    1.12,    1.12,    1.12,
  1.27,    1.27,    1.27,    1.27,
  1.87,    1.87,    1.87,    1.87,
  1.85,    1.85,    1.85,    1.85,
  1.77,    1.77,    1.77,    1.77,
  2.11,    2.11,    2.11,    2.11,
  2.41,    2.41,    2.41,    2.41,
  2.56,    2.56,    2.56,    2.56,
  1.93,    1.93,    1.93,    1.93,
  1.87,    1.87,    1.87,    1.87,
  2.149,   2.149,   2.149,   2.149,
  2.227,   2.227,   2.227,   2.227,
  2.323,   2.323,   2.323,   2.323,
  2.009,   2.009,   2.009,   2.009,
  1.975,   1.975,   1.975,   1.975,
  2.023,   2.023,   2.023,   2.023,
  1.931,   1.931,   1.931,   1.931,
  2.049,   2.049,   2.049,   2.049,
  1.991,   1.991,   1.991,   1.991,
  2.01,    2.01,    2.01,    2.01,
  2.14,    2.14,    2.14,    2.14,
  2.087,   2.087,   2.087,   2.087,
  1.921,   1.921,   1.921,   1.921,
  2.206,   2.206,   2.206,   2.206,
  2.316,   2.316,   2.316,   2.316,
  2.38,    2.38,    2.38,    2.38,
  2.467,   2.467,   2.467,   2.467,
  2.608,   2.608,   2.608,   2.608,
  2.442,   2.442,   2.442,   2.442,
  2.425,   2.425,   2.425,   2.425,
  2.66,    2.66,    2.66,    2.66,
  2.829,   2.829,   2.829,   2.829,
  2.687,   2.687,   2.687,   2.687,
  2.873,   2.873,   2.873,   2.873,
  2.695,   2.695,   2.695,   2.695,
  2.834,   2.834,   2.834,   2.834,
  2.864,   2.864,   2.864,   2.864,
  3.162,   3.162,   3.162,   3.162,
  3.11,    3.11,    3.11,    3.11,
  3.078,   3.078,   3.078,   3.078,
  3.024,   3.024,   3.024,   3.024,
  2.742,   2.742,   2.742,   2.742,
  2.639,   2.639,   2.639,   2.639,
  2.505,   2.505,   2.505,   2.505,
  2.639,   2.639,   2.639,   2.639,
  2.705,   2.705,   2.705,   2.705,
  2.825,   2.825,   2.825,   2.825,
  2.757,   2.757,   2.757,   2.757,
  2.244,   2.244,   2.244,   2.244,
  1.854,   1.854,   1.854,   1.854,
  1.874,   1.874,   1.874,   1.874,
  2.037,   2.037,   2.037,   2.037,
  2.189,   2.189,   2.189,   2.189,
  2.099,   2.099,   2.099,   2.099,
  2.247,   2.247,   2.247,   2.247,
  2.377,   2.377,   2.377,   2.377,
  2.064,   2.064,   2.064,   2.064,
  2.133,   2.133,   2.133,   2.133,
  2.149,   2.149,   2.149,   2.149,
  2.227,   2.227,   2.227,   2.227,
  2.323,   2.323,   2.323,   2.323,
  2.009,   2.009,   2.009,   2.009,
  1.975,   1.975,   1.975,   1.975,
  2.023,   2.023,   2.023,   2.023,
  1.931,   1.931,   1.931,   1.931,
  2.049,   2.049,   2.049,   2.049,
  1.991,   1.991,   1.991,   1.991,
  2.01,    2.01,    2.01,    2.01,
  2.14,    2.14,    2.14,    2.14,
  2.087,   2.087,   2.087,   2.087,
  1.921,   1.921,   1.921,   1.921,
  2.206,   2.206,   2.206,   2.206,
  2.316,   2.316,   2.316,   2.316,
  2.38,    2.38,    2.38,    2.38,
  2.467,   2.467,   2.467,   2.467,
  2.608,   2.608,   2.608,   2.608,
  2.442,   2.442,   2.442,   2.442,
  2.425,   2.425,   2.425,   2.425,
  2.66,    2.66,    2.66,    2.66,
  2.829,   2.829,   2.829,   2.829,
  2.687,   2.687,   2.687,   2.687,
  2.873,   2.873,   2.873,   2.873,
  2.695,   2.695,   2.695,   2.695,
  2.834,   2.834,   2.834,   2.834,
  2.864,   2.864,   2.864,   2.864,
  3.162,   3.162,   3.162,   3.162,
  3.11,    3.11,    3.11,    3.11,
  3.078,   3.078,   3.078,   3.078,
  3.024,   3.024,   3.024,   3.024,
  2.742,   2.742,   2.742,   2.742,
  2.639,   2.639,   2.639,   2.639,
  2.505,   2.505,   2.505,   2.505,
  2.639,   2.639,   2.639,   2.639,
  2.705,   2.705,   2.705,   2.705,
  2.825,   2.825,   2.825,   2.825,
  2.757,   2.757,   2.757,   2.757,
  2.244,   2.244,   2.244,   2.244,
  1.854,   1.854,   1.854,   1.854,
  1.874,   1.874,   1.874,   1.874,
  2.037,   2.037,   2.037,   2.037,
  2.189,   2.189,   2.189,   2.189,
  2.099,   2.099,   2.099,   2.099,
  2.247,   2.247,   2.247,   2.247,
  2.377,   2.377,   2.377,   2.377,
  2.064,   2.064,   2.064,   2.064,
  2.133,   2.133,   2.133,   2.133,
  2.149,   2.149,   2.149,   2.149,
  2.227,   2.227,   2.227,   2.227,
  2.323,   2.323,   2.323,   2.323,
  2.009,   2.009,   2.009,   2.009,
  1.975,   1.975,   1.975,   1.975,
  2.023,   2.023,   2.023,   2.023,
  1.931,   1.931,   1.931,   1.931,
  2.049,   2.049,   2.049,   2.049,
  1.991,   1.991,   1.991,   1.991,
  2.01,    2.01,    2.01,    2.01,
  2.14,    2.14,    2.14,    2.14,
  2.087,   2.087,   2.087,   2.087,
  1.921,   1.921,   1.921,   1.921,
  2.206,   2.206,   2.206,   2.206,
  2.316,   2.316,   2.316,   2.316,
  2.38,    2.38,    2.38,    2.38,
  2.467,   2.467,   2.467,   2.467,
  2.608,   2.608,   2.608,   2.608,
  2.442,   2.442,   2.442,   2.442,
  2.425,   2.425,   2.425,   2.425,
  2.66,    2.66,    2.66,    2.66,
  2.829,   2.829,   2.829,   2.829,
  2.687,   2.687,   2.687,   2.687,
  2.873,   2.873,   2.873,   2.873,
  2.695,   2.695,   2.695,   2.695,
  2.834,   2.834,   2.834,   2.834,
  2.864,   2.864,   2.864,   2.864,
  3.162,   3.162,   3.162,   3.162,
  3.11,    3.11,    3.11,    3.11,
  3.078,   3.078,   3.078,   3.078,
  3.024,   3.024,   3.024,   3.024,
  2.742,   2.742,   2.742,   2.742,
  2.639,   2.639,   2.639,   2.639,
  2.505,   2.505,   2.505,   2.505,
  2.639,   2.639,   2.639,   2.639,
  2.705,   2.705,   2.705,   2.705,
  2.825,   2.825,   2.825,   2.825,
  2.757,   2.757,   2.757,   2.757,
  2.244,   2.244,   2.244,   2.244,
  1.854,   1.854,   1.854,   1.854,
  1.874,   1.874,   1.874,   1.874,
  2.037,   2.037,   2.037,   2.037,
  2.189,   2.189,   2.189,   2.189,
  2.099,   2.099,   2.099,   2.099,
  2.247,   2.247,   2.247,   2.247,
  2.377,   2.377,   2.377,   2.377,
  2.064,   2.064,   2.064,   2.064,
  2.133,   2.133,   2.133,   2.133,
  2.149,   2.149,   2.149,   2.149,
  2.227,   2.227,   2.227,   2.227,
  2.323,   2.323,   2.323,   2.323,
  2.009,   2.009,   2.009,   2.009,
  1.975,   1.975,   1.975,   1.975,
  2.023,   2.023,   2.023,   2.023,
  1.931,   1.931,   1.931,   1.931,
  2.049,   2.049,   2.049,   2.049,
  1.991,   1.991,   1.991,   1.991,
  2.01,    2.01,    2.01,    2.01,
  2.14,    2.14,    2.14,    2.14,
  2.087,   2.087,   2.087,   2.087,
  1.921,   1.921,   1.921,   1.921,
  2.206,   2.206,   2.206,   2.206,
  2.316,   2.316,   2.316,   2.316,
  2.38,    2.38,    2.38,    2.38,
  2.467,   2.467,   2.467,   2.467,
  2.608,   2.608,   2.608,   2.608,
  2.442,   2.442,   2.442,   2.442,
  2.425,   2.425,   2.425,   2.425,
  2.66,    2.66,    2.66,    2.66,
  2.829,   2.829,   2.829,   2.829,
  2.687,   2.687,   2.687,   2.687,
  2.873,   2.873,   2.873,   2.873,
  2.695,   2.695,   2.695,   2.695,
  2.834,   2.834,   2.834,   2.834,
  2.864,   2.864,   2.864,   2.864,
  3.162,   3.162,   3.162,   3.162,
  3.11,    3.11,    3.11,    3.11,
  3.078,   3.078,   3.078,   3.078,
  3.024,   3.024,   3.024,   3.024,
  3.01,    3.01,    3.01,    3.01,
  2.79,    2.79,    2.79,    2.79,
  2.52,    2.52,    2.52,    2.52,
  2.15,    2.15,    2.15,    2.15,
  1.9,     1.9,     1.9,     1.9,
  1.77,    1.77,    1.77,    1.77,
  1.99,    1.99,    1.99,    1.99,
  2.14,    2.14,    2.14,    2.14,
  1.42,    1.42,    1.42,    1.42,
  1.36,    1.36,    1.36,    1.36,
  1.85,    1.85,    1.85,    1.85,
  1.71,    1.71,    1.71,    1.71,
  1.82,    1.82,    1.82,    1.82,
  2.09,    2.09,    2.09,    2.09,
  2.16,    2.16,    2.16,    2.16,
  2.1,     2.1,     2.1,     2.1,
  1.8,     1.8,     1.8,     1.8,
  1.81,    1.81,    1.81,    1.81,
  1.9,     1.9,     1.9,     1.9,
  2.26,    2.26,    2.26,    2.26,
  0.54,    0.54,    0.54,    0.54,
  0.22,    0.22,    0.22,    0.22,
  0.95,    0.95,    0.95,    0.95,
  0.2,     0.2,     0.2,     0.2,
  0.91,    0.91,    0.91,    0.91,
  0.55,    0.55,    0.55,    0.55,
  0.75,    0.75,    0.75,    0.75,
  1.39,    1.39,    1.39,    1.39,
  1.11,    1.11,    1.11,    1.11,
  0.45,    0.45,    0.45,    0.45,
  0.58,    0.58,    0.58,    0.58,
  0.64,    0.64,    0.64,    0.64,
  1.24,    1.24,    1.24,    1.24,
  1.65,    1.65,    1.65,    1.65,
  1.96,    1.96,    1.96,    1.96,
  2.21,    2.21,    2.21,    2.21,
  1.77,    1.77,    1.77,    1.77,
  2.32,    2.32,    2.32,    2.32,
  2.57,    2.57,    2.57,    2.57,
  2.85,    2.85,    2.85,    2.85,
  2.96,    2.96,    2.96,    2.96,
  2.29,    2.29,    2.29,    2.29,
  2.81,    2.81,    2.81,    2.81,
  2.73,    2.73,    2.73,    2.73,
  2.28,    2.28,    2.28,    2.28,
  2.81,    2.81,    2.81,    2.81,
  3.12,    3.12,    3.12,    3.12,
  2.65,    2.65,    2.65,    2.65,
  2.32,    2.32,    2.32,    2.32,
  2.76,    2.76,    2.76,    2.76,
  1.4,     1.4,     1.4,     1.4,
  1.65,    1.65,    1.65,    1.65,
  2.11,    2.11,    2.11,    2.11,
  2,       2,       2,       2,
  2.32,    2.32,    2.32,    2.32,
  1.97,    1.97,    1.97,    1.97,
  1.46,    1.46,    1.46,    1.46,
  1.26,    1.26,    1.26,    1.26,
  1.9,     1.9,     1.9,     1.9,
  1.65,    1.65,    1.65,    1.65,
  1.42,    1.42,    1.42,    1.42,
  1.82,    1.82,    1.82,    1.82,
  1.41,    1.41,    1.41,    1.41,
  0.55,    0.55,    0.55,    0.55,
  0.97,    0.97,    0.97,    0.97,
  1.1,     1.1,     1.1,     1.1,
  1.23,    1.23,    1.23,    1.23,
  1.63,    1.63,    1.63,    1.63,
  2.02,    2.02,    2.02,    2.02,
  1.74,    1.74,    1.74,    1.74,
  1.49,    1.49,    1.49,    1.49,
  1.46,    1.46,    1.46,    1.46,
  1.18,    1.18,    1.18,    1.18,
  1.55,    1.55,    1.55,    1.55,
  1.64,    1.64,    1.64,    1.64,
  1.45,    1.45,    1.45,    1.45,
  1.75,    1.75,    1.75,    1.75,
  2.11,    2.11,    2.11,    2.11,
  2.9,     2.9,     2.9,     2.9,
  3.31,    3.31,    3.31,    3.31,
  2.98,    2.98,    2.98,    2.98,
  3.17,    3.17,    3.17,    3.17,
  3.45,    3.45,    3.45,    3.45,
  3.44,    3.44,    3.44,    3.44,
  2.99,    2.99,    2.99,    2.99,
  3.31,    3.31,    3.31,    3.31,
  3.22,    3.22,    3.22,    3.22,
  3.53,    3.53,    3.53,    3.53,
  3.24,    3.24,    3.24,    3.24,
  3.3,     3.3,     3.3,     3.3,
  2.82,    2.82,    2.82,    2.82,
  3.02,    3.02,    3.02,    3.02,
  3.17,    3.17,    3.17,    3.17,
  3.18,    3.18,    3.18,    3.18,
  2.97,    2.97,    2.97,    2.97,
  2.59,    2.59,    2.59,    2.59,
  2.64,    2.64,    2.64,    2.64,
  1.75,    1.75,    1.75,    1.75,
  1.73,    1.73,    1.73,    1.73,
  3.27,    3.27,    3.27,    3.27,
  3.06,    3.06,    3.06,    3.06,
  3.34,    3.34,    3.34,    3.34,
  3.33,    3.33,    3.33,    3.33,
  3.24,    3.24,    3.24,    3.24,
  3.15,    3.15,    3.15,    3.15,
  3.73,    3.73,    3.73,    3.73,
  3.31,    3.31,    3.31,    3.31,
  2.94,    2.94,    2.94,    2.94,
  2.09,    2.09,    2.09,    2.09,
  2.26,    2.26,    2.26,    2.26,
  2.57,    2.57,    2.57,    2.57,
  2.54,    2.54,    2.54,    2.54,
  2.65,    2.65,    2.65,    2.65,
  2.84,    2.84,    2.84,    2.84,
  2.55,    2.55,    2.55,    2.55,
  2.86,    2.86,    2.86,    2.86,
  2.52,    2.52,    2.52,    2.52,
  2.59,    2.59,    2.59,    2.59,
  2.27,    2.27,    2.27,    2.27,
  2.38,    2.38,    2.38,    2.38,
  2.26,    2.26,    2.26,    2.26,
  2.85,    2.85,    2.85,    2.85,
  2.3,     2.3,     2.3,     2.3,
  2.28,    2.28,    2.28,    2.28,
  2.71,    2.71,    2.71,    2.71,
  2.5,     2.5,     2.5,     2.5,
  2.74,    2.74,    2.74,    2.74,
  2.98,    2.98,    2.98,    2.98,
  2.87,    2.87,    2.87,    2.87,
  2.37,    2.37,    2.37,    2.37,
  3.1,     3.1,     3.1,     3.1,
  2.87,    2.87,    2.87,    2.87,
  2.91,    2.91,    2.91,    2.91,
  3.02,    3.02,    3.02,    3.02,
  2.87,    2.87,    2.87,    2.87,
  2.6,     2.6,     2.6,     2.6,
  3.53,    3.53,    3.53,    3.53,
  3.53,    3.53,    3.53,    3.53,
  3.4,     3.4,     3.4,     3.4,
  2.87,    2.87,    2.87,    2.87,
  3.62,    3.62,    3.62,    3.62,
  3.33,    3.33,    3.33,    3.33,
  3.56,    3.56,    3.56,    3.56,
  3.78,    3.78,    3.78,    3.78,
  3.67,    3.67,    3.67,    3.67,
  2.99,    2.99,    2.99,    2.99,
  3.19,    3.19,    3.19,    3.19,
  2.7,     2.7,     2.7,     2.7,
  1.69,    1.69,    1.69,    1.69,
  2.53,    2.53,    2.53,    2.53,
  2.42,    2.42,    2.42,    2.42,
  2.05,    2.05,    2.05,    2.05,
  1.43,    1.43,    1.43,    1.43,
  1.03,    1.03,    1.03,    1.03,
  1.07,    1.07,    1.07,    1.07,
  1.59,    1.59,    1.59,    1.59,
  1.75,    1.75,    1.75,    1.75,
  0.98,    0.98,    0.98,    0.98,
  1.83,    1.83,    1.83,    1.83,
  1.72,    1.72,    1.72,    1.72,
  1.41,    1.41,    1.41,    1.41,
  1.17,    1.17,    1.17,    1.17,
  0.65,    0.65,    0.65,    0.65,
  0.71,    0.71,    0.71,    0.71,
  0.39,    0.39,    0.39,    0.39,
  0.43,    0.43,    0.43,    0.43,
  0.72,    0.72,    0.72,    0.72,
  0.5,     0.5,     0.5,     0.5,
  0.46,    0.46,    0.46,    0.46,
  0.76,    0.76,    0.76,    0.76,
  0.97,    0.97,    0.97,    0.97,
  1.02,    1.02,    1.02,    1.02,
  0.63,    0.63,    0.63,    0.63,
  0.44,    0.44,    0.44,    0.44,
  0.73,    0.73,    0.73,    0.73,
  0.98,    0.98,    0.98,    0.98,
  1.09,    1.09,    1.09,    1.09,
  1.52,    1.52,    1.52,    1.52,
  0.95,    0.95,    0.95,    0.95,
  1.29,    1.29,    1.29,    1.29,
  1.78,    1.78,    1.78,    1.78,
  2.02,    2.02,    2.02,    2.02,
  2.13,    2.13,    2.13,    2.13,
  1.44,    1.44,    1.44,    1.44,
  1.33,    1.33,    1.33,    1.33,
  1.73,    1.73,    1.73,    1.73,
  2.42,    2.42,    2.42,    2.42,
  1.53,    1.53,    1.53,    1.53,
  2.99,    2.99,    2.99,    2.99,
  2.88,    2.88,    2.88,    2.88,
  2.73,    2.73,    2.73,    2.73,
  1.71,    1.71,    1.71,    1.71,
  2.39,    2.39,    2.39,    2.39,
  2.25,    2.25,    2.25,    2.25,
  2.35,    2.35,    2.35,    2.35,
  2.51,    2.51,    2.51,    2.51,
  2.58,    2.58,    2.58,    2.58,
  3.09,    3.09,    3.09,    3.09,
  3.08,    3.08,    3.08,    3.08,
  2.73,    2.73,    2.73,    2.73,
  1.94,    1.94,    1.94,    1.94,
  1.87,    1.87,    1.87,    1.87,
  2.3,     2.3,     2.3,     2.3,
  2.67,    2.67,    2.67,    2.67,
  2.61,    2.61,    2.61,    2.61,
  2.7,     2.7,     2.7,     2.7,
  2.83,    2.83,    2.83,    2.83,
  2.45,    2.45,    2.45,    2.45,
  2.38,    2.38,    2.38,    2.38,
  2.67,    2.67,    2.67,    2.67,
  2.76,    2.76,    2.76,    2.76,
  2.35,    2.35,    2.35,    2.35,
  2.25,    2.25,    2.25,    2.25,
  1.93,    1.93,    1.93,    1.93,
  2.07,    2.07,    2.07,    2.07,
  2.08,    2.08,    2.08,    2.08,
  2.08,    2.08,    2.08,    2.08,
  1.59,    1.59,    1.59,    1.59,
  1.87,    1.87,    1.87,    1.87,
  2.08,    2.08,    2.08,    2.08,
  2.31,    2.31,    2.31,    2.31,
  2.73,    2.73,    2.73,    2.73,
  3.29,    3.29,    3.29,    3.29,
  3.16,    3.16,    3.16,    3.16,
  3.75,    3.75,    3.75,    3.75,
  3.09,    3.09,    3.09,    3.09,
  3.11,    3.11,    3.11,    3.11,
  2.27,    2.27,    2.27,    2.27,
  2.63,    2.63,    2.63,    2.63,
  2.57,    2.57,    2.57,    2.57,
  2.58,    2.58,    2.58,    2.58,
  2.46,    2.46,    2.46,    2.46,
  2.69,    2.69,    2.69,    2.69,
  2.31,    2.31,    2.31,    2.31,
  2.72,    2.72,    2.72,    2.72,
  2.18,    2.18,    2.18,    2.18,
  2.76,    2.76,    2.76,    2.76,
  2.7,     2.7,     2.7,     2.7,
  3.12,    3.12,    3.12,    3.12,
  3.41,    3.41,    3.41,    3.41,
  3.23,    3.23,    3.23,    3.23,
  3.36,    3.36,    3.36,    3.36,
  2.87,    2.87,    2.87,    2.87,
  3.42,    3.42,    3.42,    3.42,
  3.69,    3.69,    3.69,    3.69,
  4.12,    4.12,    4.12,    4.12,
  3.9,     3.9,     3.9,     3.9,
  3.4,     3.4,     3.4,     3.4,
  2.08,    2.08,    2.08,    2.08,
  1.94,    1.94,    1.94,    1.94,
  1.74,    1.74,    1.74,    1.74,
  2.44,    2.44,    2.44,    2.44,
  2.28,    2.28,    2.28,    2.28,
  2.19,    2.19,    2.19,    2.19,
  2.31,    2.31,    2.31,    2.31,
  1.98,    1.98,    1.98,    1.98,
  1.61,    1.61,    1.61,    1.61,
  1.76,    1.76,    1.76,    1.76,
  1.52,    1.52,    1.52,    1.52,
  1.72,    1.72,    1.72,    1.72,
  1.81,    1.81,    1.81,    1.81,
  1.69,    1.69,    1.69,    1.69,
  1.54,    1.54,    1.54,    1.54,
  0.22,    0.22,    0.22,    0.22,
  0.21,    0.21,    0.21,    0.21,
  0.51,    0.51,    0.51,    0.51,
  1.03,    1.03,    1.03,    1.03,
  0.93,    0.93,    0.93,    0.93,
  0.58,    0.58,    0.58,    0.58,
  0.62,    0.62,    0.62,    0.62,
  0.6,     0.6,     0.6,     0.6,
  0.45,    0.45,    0.45,    0.45,
  0.55,    0.55,    0.55,    0.55,
  1.57,    1.57,    1.57,    1.57,
  0.99,    0.99,    0.99,    0.99,
  1.01,    1.01,    1.01,    1.01,
  1.82,    1.82,    1.82,    1.82,
  1.65,    1.65,    1.65,    1.65,
  0.93,    0.93,    0.93,    0.93,
  1.76,    1.76,    1.76,    1.76,
  0.67,    0.67,    0.67,    0.67,
  1.17,    1.17,    1.17,    1.17,
  0.83,    0.83,    0.83,    0.83,
  1.32,    1.32,    1.32,    1.32,
  0.98,    0.98,    0.98,    0.98,
  1.07,    1.07,    1.07,    1.07,
  1.68,    1.68,    1.68,    1.68,
  2.43,    2.43,    2.43,    2.43,
  1.96,    1.96,    1.96,    1.96,
  1.76,    1.76,    1.76,    1.76,
  1.92,    1.92,    1.92,    1.92,
  1.4,     1.4,     1.4,     1.4,
  1.98,    1.98,    1.98,    1.98,
  1.21,    1.21,    1.21,    1.21,
  0.85,    0.85,    0.85,    0.85,
  1.27,    1.27,    1.27,    1.27,
  1.24,    1.24,    1.24,    1.24,
  1.58,    1.58,    1.58,    1.58,
  2.08,    2.08,    2.08,    2.08,
  2.23,    2.23,    2.23,    2.23,
  2.35,    2.35,    2.35,    2.35,
  2.4,     2.4,     2.4,     2.4,
  2.38,    2.38,    2.38,    2.38,
  2.36,    2.36,    2.36,    2.36,
  2.46,    2.46,    2.46,    2.46,
  2.44,    2.44,    2.44,    2.44,
  2.4,     2.4,     2.4,     2.4,
  2.46,    2.46,    2.46,    2.46,
  2.54,    2.54,    2.54,    2.54,
  2.53,    2.53,    2.53,    2.53,
  2.53,    2.53,    2.53,    2.53,
  2.55,    2.55,    2.55,    2.55,
  2.42,    2.42,    2.42,    2.42,
  2.48,    2.48,    2.48,    2.48,
  2.57,    2.57,    2.57,    2.57,
  2.3,     2.3,     2.3,     2.3,
  2.27,    2.27,    2.27,    2.27,
  2.27,    2.27,    2.27,    2.27,
  2.55,    2.55,    2.55,    2.55,
  3.21,    3.21,    3.21,    3.21,
  3.07,    3.07,    3.07,    3.07,
  3.86,    3.86,    3.86,    3.86,
  3.87,    3.87,    3.87,    3.87,
  3.98,    3.98,    3.98,    3.98,
  3.84,    3.84,    3.84,    3.84,
  3.86,    3.86,    3.86,    3.86,
  3.52,    3.52,    3.52,    3.52,
  3.85,    3.85,    3.85,    3.85,
  3.48,    3.48,    3.48,    3.48,
  2.52,    2.52,    2.52,    2.52,
  2.69,    2.69,    2.69,    2.69,
  2.82,    2.82,    2.82,    2.82,
  3.57,    3.57,    3.57,    3.57,
  2.81,    2.81,    2.81,    2.81,
  2.85,    2.85,    2.85,    2.85,
  2.82,    2.82,    2.82,    2.82,
  2.81,    2.81,    2.81,    2.81,
  2.82,    2.82,    2.82,    2.82,
  2.84,    2.84,    2.84,    2.84,
  2.9,     2.9,     2.9,     2.9,
  2.88,    2.88,    2.88,    2.88,
  2.66,    2.66,    2.66,    2.66,
  2.32,    2.32,    2.32,    2.32,
  1.85,    1.85,    1.85,    1.85,
  2.29,    2.29,    2.29,    2.29,
  2.25,    2.25,    2.25,    2.25,
  2.2,     2.2,     2.2,     2.2,
  2.48,    2.48,    2.48,    2.48,
  1.43,    1.43,    1.43,    1.43,
  1.15,    1.15,    1.15,    1.15,
  2.2,     2.2,     2.2,     2.2,
  2.68,    2.68,    2.68,    2.68,
  2.35,    2.35,    2.35,    2.35,
  2.22,    2.22,    2.22,    2.22,
  2.13,    2.13,    2.13,    2.13,
  1.56,    1.56,    1.56,    1.56,
  1.25,    1.25,    1.25,    1.25,
  1.68,    1.68,    1.68,    1.68,
  1.79,    1.79,    1.79,    1.79,
  2.9,     2.9,     2.9,     2.9,
  2.01,    2.01,    2.01,    2.01,
  2.48,    2.48,    2.48,    2.48,
  2.84,    2.84,    2.84,    2.84,
  2.1,     2.1,     2.1,     2.1,
  2.38,    2.38,    2.38,    2.38,
  2.45,    2.45,    2.45,    2.45,
  2.11,    2.11,    2.11,    2.11,
  2.68,    2.68,    2.68,    2.68,
  2.95,    2.95,    2.95,    2.95,
  2.69,    2.69,    2.69,    2.69,
  3.36,    3.36,    3.36,    3.36,
  3.62,    3.62,    3.62,    3.62,
  4.13,    4.13,    4.13,    4.13,
  4.28,    4.28,    4.28,    4.28,
  3.98,    3.98,    3.98,    3.98,
  3.81,    3.81,    3.81,    3.81,
  3.9,     3.9,     3.9,     3.9,
  3.86,    3.86,    3.86,    3.86,
  3.55,    3.55,    3.55,    3.55,
  3.08,    3.08,    3.08,    3.08,
  3.73,    3.73,    3.73,    3.73,
  3.22,    3.22,    3.22,    3.22,
  3.93,    3.93,    3.93,    3.93,
  4.08,    4.08,    4.08,    4.08,
  4.08,    4.08,    4.08,    4.08,
  4.4,     4.4,     4.4,     4.4,
  3.37,    3.37,    3.37,    3.37,
  2.67,    2.67,    2.67,    2.67,
  1.52,    1.52,    1.52,    1.52,
  1.99,    1.99,    1.99,    1.99,
  1.38,    1.38,    1.38,    1.38,
  1.59,    1.59,    1.59,    1.59,
  1.9,     1.9,     1.9,     1.9,
  2.44,    2.44,    2.44,    2.44,
  3.48,    3.48,    3.48,    3.48,
  2.38,    2.38,    2.38,    2.38,
  2.12,    2.12,    2.12,    2.12,
  2.56,    2.56,    2.56,    2.56,
  2.92,    2.92,    2.92,    2.92,
  2.72,    2.72,    2.72,    2.72,
  3.56,    3.56,    3.56,    3.56,
  4.09,    4.09,    4.09,    4.09,
  3.49,    3.49,    3.49,    3.49,
  3.81,    3.81,    3.81,    3.81,
  3.35,    3.35,    3.35,    3.35,
  2.83,    2.83,    2.83,    2.83,
  3.13,    3.13,    3.13,    3.13,
  2.9,     2.9,     2.9,     2.9,
  2.94,    2.94,    2.94,    2.94,
  2.44,    2.44,    2.44,    2.44,
  2.62,    2.62,    2.62,    2.62,
  3.42,    3.42,    3.42,    3.42,
  3.28,    3.28,    3.28,    3.28,
  3.57,    3.57,    3.57,    3.57,
  3.33,    3.33,    3.33,    3.33,
  3.61,    3.61,    3.61,    3.61,
  4,       4,       4,       4,
  4.25,    4.25,    4.25,    4.25,
  3.91,    3.91,    3.91,    3.91,
  4.24,    4.24,    4.24,    4.24,
  3.7,     3.7,     3.7,     3.7,
  5.19,    5.19,    5.19,    5.19,
  4.17,    4.17,    4.17,    4.17,
  5.06,    5.06,    5.06,    5.06,
  5.15,    5.15,    5.15,    5.15,
  4.84,    4.84,    4.84,    4.84,
  3.18,    3.18,    3.18,    3.18,
  3.73,    3.73,    3.73,    3.73,
  4.24,    4.24,    4.24,    4.24,
  4.18,    4.18,    4.18,    4.18,
  3.37,    3.37,    3.37,    3.37,
  3.53,    3.53,    3.53,    3.53,
  3.83,    3.83,    3.83,    3.83,
  3.57,    3.57,    3.57,    3.57,
  3.62,    3.62,    3.62,    3.62,
  2.71,    2.71,    2.71,    2.71,
  2.79,    2.79,    2.79,    2.79,
  1.87,    1.87,    1.87,    1.87,
  1.02,    1.02,    1.02,    1.02,
  2.31,    2.31,    2.31,    2.31,
  3.78,    3.78,    3.78,    3.78,
  2.64,    2.64,    2.64,    2.64,
  2.37,    2.37,    2.37,    2.37,
  1.89,    1.89,    1.89,    1.89,
  1.87,    1.87,    1.87,    1.87,
  2.2,     2.2,     2.2,     2.2,
  2.65,    2.65,    2.65,    2.65,
  2.78,    2.78,    2.78,    2.78,
  2.85,    2.85,    2.85,    2.85,
  2.36,    2.36,    2.36,    2.36,
  2.14,    2.14,    2.14,    2.14,
  1.92,    1.92,    1.92,    1.92,
  2.01,    2.01,    2.01,    2.01,
  2.03,    2.03,    2.03,    2.03,
  2.41,    2.41,    2.41,    2.41,
  2.42,    2.42,    2.42,    2.42,
  2.43,    2.43,    2.43,    2.43,
  2.49,    2.49,    2.49,    2.49,
  2.69,    2.69,    2.69,    2.69,
  2.84,    2.84,    2.84,    2.84,
  3.04,    3.04,    3.04,    3.04,
  3.51,    3.51,    3.51,    3.51,
  3.4,     3.4,     3.4,     3.4,
  4.11,    4.11,    4.11,    4.11,
  4.36,    4.36,    4.36,    4.36,
  4.93,    4.93,    4.93,    4.93,
  5.46,    5.46,    5.46,    5.46,
  4.96,    4.96,    4.96,    4.96,
  5.64,    5.64,    5.64,    5.64,
  5.58,    5.58,    5.58,    5.58,
  5.51,    5.51,    5.51,    5.51,
  4.9,     4.9,     4.9,     4.9,
  5.73,    5.73,    5.73,    5.73,
  4.87,    4.87,    4.87,    4.87,
  4.59,    4.59,    4.59,    4.59,
  4.59,    4.59,    4.59,    4.59,
  4.24,    4.24,    4.24,    4.24,
  4.66,    4.66,    4.66,    4.66,
  4.6,     4.6,     4.6,     4.6,
  4,       4,       4,       4,
  4.05,    4.05,    4.05,    4.05,
  3.18,    3.18,    3.18,    3.18,
  3.86,    3.86,    3.86,    3.86,
  3.31,    3.31,    3.31,    3.31,
  3.93,    3.93,    3.93,    3.93,
  3.57,    3.57,    3.57,    3.57,
  3.25,    3.25,    3.25,    3.25,
  3.06,    3.06,    3.06,    3.06,
  2.8,     2.8,     2.8,     2.8,
  2.6,     2.6,     2.6,     2.6,
  2.57,    2.57,    2.57,    2.57,
  2.18,    2.18,    2.18,    2.18,
  2.27,    2.27,    2.27,    2.27,
  2.39,    2.39,    2.39,    2.39,
  2.06,    2.06,    2.06,    2.06,
  1.88,    1.88,    1.88,    1.88,
  1.71,    1.71,    1.71,    1.71,
  1.89,    1.89,    1.89,    1.89,
  2.2,     2.2,     2.2,     2.2,
  1.75,    1.75,    1.75,    1.75,
  1.8,     1.8,     1.8,     1.8,
  1.64,    1.64,    1.64,    1.64,
  1.71,    1.71,    1.71,    1.71,
  1.94,    1.94,    1.94,    1.94,
  1.94,    1.94,    1.94,    1.94,
  2.14,    2.14,    2.14,    2.14,
  2.24,    2.24,    2.24,    2.24,
  2.13,    2.13,    2.13,    2.13,
  2.48,    2.48,    2.48,    2.48,
  2.27,    2.27,    2.27,    2.27,
  2.85,    2.85,    2.85,    2.85,
  3.72,    3.72,    3.72,    3.72,
  3.37,    3.37,    3.37,    3.37,
  3.65,    3.65,    3.65,    3.65,
  3.22,    3.22,    3.22,    3.22,
  2.7,     2.7,     2.7,     2.7,
  2.78,    2.78,    2.78,    2.78,
  3.88,    3.88,    3.88,    3.88,
  3.98,    3.98,    3.98,    3.98,
  4.33,    4.33,    4.33,    4.33,
  4.46,    4.46,    4.46,    4.46,
  3.88,    3.88,    3.88,    3.88,
  4.89,    4.89,    4.89,    4.89,
  4.43,    4.43,    4.43,    4.43,
  4.95,    4.95,    4.95,    4.95,
  5.44,    5.44,    5.44,    5.44,
  5.34,    5.34,    5.34,    5.34,
  4.61,    4.61,    4.61,    4.61,
  4.93,    4.93,    4.93,    4.93,
  4.85,    4.85,    4.85,    4.85,
  4.85,    4.85,    4.85,    4.85,
  4.95,    4.95,    4.95,    4.95,
  4.22,    4.22,    4.22,    4.22,
  4.92,    4.92,    4.92,    4.92,
  4.7,     4.7,     4.7,     4.7,
  3.93,    3.93,    3.93,    3.93,
  3.7,     3.7,     3.7,     3.7,
  3.71,    3.71,    3.71,    3.71,
  3.44,    3.44,    3.44,    3.44,
  3.38,    3.38,    3.38,    3.38,
  3.69,    3.69,    3.69,    3.69,
  3.21,    3.21,    3.21,    3.21,
  3.4,     3.4,     3.4,     3.4,
  2.97,    2.97,    2.97,    2.97,
  3.2,     3.2,     3.2,     3.2,
  3.1,     3.1,     3.1,     3.1,
  3.3,     3.3,     3.3,     3.3,
  3.32,    3.32,    3.32,    3.32,
  3.19,    3.19,    3.19,    3.19,
  3.07,    3.07,    3.07,    3.07,
  3.27,    3.27,    3.27,    3.27,
  2.9,     2.9,     2.9,     2.9,
  3.51,    3.51,    3.51,    3.51,
  2.73,    2.73,    2.73,    2.73,
  2.66,    2.66,    2.66,    2.66,
  2.9,     2.9,     2.9,     2.9,
  3.09,    3.09,    3.09,    3.09,
  2.76,    2.76,    2.76,    2.76,
  3.14,    3.14,    3.14,    3.14,
  3.47,    3.47,    3.47,    3.47,
  3.77,    3.77,    3.77,    3.77,
  4.4,     4.4,     4.4,     4.4,
  4.72,    4.72,    4.72,    4.72,
  4,       4,       4,       4,
  3.94,    3.94,    3.94,    3.94,
  4.45,    4.45,    4.45,    4.45,
  3.95,    3.95,    3.95,    3.95,
  4.22,    4.22,    4.22,    4.22,
  4.47,    4.47,    4.47,    4.47,
  3.76,    3.76,    3.76,    3.76,
  4.02,    4.02,    4.02,    4.02,
  4.33,    4.33,    4.33,    4.33,
  5.1,     5.1,     5.1,     5.1,
  4.52,    4.52,    4.52,    4.52,
  4.46,    4.46,    4.46,    4.46,
  4.21,    4.21,    4.21,    4.21,
  4.22,    4.22,    4.22,    4.22,
  4.4,     4.4,     4.4,     4.4,
  3.76,    3.76,    3.76,    3.76,
  3.63,    3.63,    3.63,    3.63,
  3.78,    3.78,    3.78,    3.78,
  2.97,    2.97,    2.97,    2.97,
  2.86,    2.86,    2.86,    2.86,
  1.92,    1.92,    1.92,    1.92,
  2.83,    2.83,    2.83,    2.83,
  2.22,    2.22,    2.22,    2.22,
  1.9,     1.9,     1.9,     1.9,
  1.98,    1.98,    1.98,    1.98,
  1.66,    1.66,    1.66,    1.66,
  1.82,    1.82,    1.82,    1.82,
  2.31,    2.31,    2.31,    2.31,
  2.24,    2.24,    2.24,    2.24,
  2.13,    2.13,    2.13,    2.13,
  2.26,    2.26,    2.26,    2.26,
  2.23,    2.23,    2.23,    2.23,
  2.18,    2.18,    2.18,    2.18,
  2.36,    2.36,    2.36,    2.36,
  2.15,    2.15,    2.15,    2.15,
  1.91,    1.91,    1.91,    1.91,
  1.79,    1.79,    1.79,    1.79,
  2.06,    2.06,    2.06,    2.06,
  1.83,    1.83,    1.83,    1.83,
  1.88,    1.88,    1.88,    1.88,
  1.82,    1.82,    1.82,    1.82,
  1.51,    1.51,    1.51,    1.51,
  1.44,    1.44,    1.44,    1.44,
  1.86,    1.86,    1.86,    1.86,
  2.78,    2.78,    2.78,    2.78,
  3.22,    3.22,    3.22,    3.22,
  3.96,    3.96,    3.96,    3.96,
  3.38,    3.38,    3.38,    3.38,
  3.93,    3.93,    3.93,    3.93,
  3.49,    3.49,    3.49,    3.49,
  4,       4,       4,       4,
  3.96,    3.96,    3.96,    3.96,
  4.32,    4.32,    4.32,    4.32,
  3.82,    3.82,    3.82,    3.82,
  3.8,     3.8,     3.8,     3.8,
  3.67,    3.67,    3.67,    3.67,
  3.5,     3.5,     3.5,     3.5,
  3.31,    3.31,    3.31,    3.31,
  3.27,    3.27,    3.27,    3.27,
  2.96,    2.96,    2.96,    2.96,
  2.22,    2.22,    2.22,    2.22,
  1.96,    1.96,    1.96,    1.96,
  1.92,    1.92,    1.92,    1.92,
  2.36,    2.36,    2.36,    2.36,
  1.71,    1.71,    1.71,    1.71,
  1.27,    1.27,    1.27,    1.27,
  0.78,    0.78,    0.78,    0.78,
  1.16,    1.16,    1.16,    1.16,
  1.37,    1.37,    1.37,    1.37,
  1.42,    1.42,    1.42,    1.42,
  1.49,    1.49,    1.49,    1.49,
  1.78,    1.78,    1.78,    1.78,
  1.72,    1.72,    1.72,    1.72,
  2.03,    2.03,    2.03,    2.03,
  2.24,    2.24,    2.24,    2.24,
  2.77,    2.77,    2.77,    2.77,
  2.76,    2.76,    2.76,    2.76,
  2.74,    2.74,    2.74,    2.74,
  2.94,    2.94,    2.94,    2.94,
  2.73,    2.73,    2.73,    2.73,
  2.68,    2.68,    2.68,    2.68,
  2.04,    2.04,    2.04,    2.04,
  1.99,    1.99,    1.99,    1.99,
  2.68,    2.68,    2.68,    2.68,
  2.75,    2.75,    2.75,    2.75,
  2.63,    2.63,    2.63,    2.63,
  2.35,    2.35,    2.35,    2.35,
  2.23,    2.23,    2.23,    2.23,
  2.12,    2.12,    2.12,    2.12,
  2.25,    2.25,    2.25,    2.25,
  2.42,    2.42,    2.42,    2.42,
  2.42,    2.42,    2.42,    2.42,
  2.47,    2.47,    2.47,    2.47,
  2.71,    2.71,    2.71,    2.71,
  2.67,    2.67,    2.67,    2.67,
  2.83,    2.83,    2.83,    2.83,
  2.98,    2.98,    2.98,    2.98,
  2.7,     2.7,     2.7,     2.7,
  2.64,    2.64,    2.64,    2.64,
  2.62,    2.62,    2.62,    2.62,
  2.47,    2.47,    2.47,    2.47,
  2.87,    2.87,    2.87,    2.87,
  3.54,    3.54,    3.54,    3.54,
  3.41,    3.41,    3.41,    3.41,
  2.96,    2.96,    2.96,    2.96,
  2.07,    2.07,    2.07,    2.07,
  1.45,    1.45,    1.45,    1.45,
  1.4,     1.4,     1.4,     1.4,
  1.24,    1.24,    1.24,    1.24,
  1.78,    1.78,    1.78,    1.78,
  1.09,    1.09,    1.09,    1.09,
  1.16,    1.16,    1.16,    1.16,
  1.49,    1.49,    1.49,    1.49,
  1.45,    1.45,    1.45,    1.45,
  1.4,     1.4,     1.4,     1.4,
  1.35,    1.35,    1.35,    1.35,
  1.79,    1.79,    1.79,    1.79,
  1.73,    1.73,    1.73,    1.73,
  2.1,     2.1,     2.1,     2.1,
  2.02,    2.02,    2.02,    2.02,
  2.03,    2.03,    2.03,    2.03,
  1.96,    1.96,    1.96,    1.96,
  2.03,    2.03,    2.03,    2.03,
  1.87,    1.87,    1.87,    1.87,
  2.23,    2.23,    2.23,    2.23,
  2.12,    2.12,    2.12,    2.12,
  2.21,    2.21,    2.21,    2.21,
  2.31,    2.31,    2.31,    2.31,
  2.45,    2.45,    2.45,    2.45,
  2.58,    2.58,    2.58,    2.58,
  2.31,    2.31,    2.31,    2.31,
  2.69,    2.69,    2.69,    2.69,
  2.42,    2.42,    2.42,    2.42,
  2.21,    2.21,    2.21,    2.21,
  1.98,    1.98,    1.98,    1.98,
  1.49,    1.49,    1.49,    1.49,
  1.6,     1.6,     1.6,     1.6,
  1.42,    1.42,    1.42,    1.42,
  1.66,    1.66,    1.66,    1.66,
  1.68,    1.68,    1.68,    1.68,
  1.25,    1.25,    1.25,    1.25,
  1.59,    1.59,    1.59,    1.59,
  1.91,    1.91,    1.91,    1.91,
  2.06,    2.06,    2.06,    2.06,
  1.86,    1.86,    1.86,    1.86,
  1.36,    1.36,    1.36,    1.36,
  1.4,     1.4,     1.4,     1.4,
  1.35,    1.35,    1.35,    1.35,
  1.2,     1.2,     1.2,     1.2,
  1.4,     1.4,     1.4,     1.4,
  2.24,    2.24,    2.24,    2.24,
  1.62,    1.62,    1.62,    1.62,
  1.11,    1.11,    1.11,    1.11,
  2.86,    2.86,    2.86,    2.86,
  3.58,    3.58,    3.58,    3.58,
  3.72,    3.72,    3.72,    3.72,
  1.65,    1.65,    1.65,    1.65,
  0.53,    0.53,    0.53,    0.53,
  0.82,    0.82,    0.82,    0.82,
  1.06,    1.06,    1.06,    1.06,
  1.57,    1.57,    1.57,    1.57,
  1.75,    1.75,    1.75,    1.75,
  1.67,    1.67,    1.67,    1.67,
  2.29,    2.29,    2.29,    2.29,
  2.22,    2.22,    2.22,    2.22,
  1.63,    1.63,    1.63,    1.63,
  2.23,    2.23,    2.23,    2.23,
  2.34,    2.34,    2.34,    2.34,
  2.44,    2.44,    2.44,    2.44,
  2.34,    2.34,    2.34,    2.34,
  2.33,    2.33,    2.33,    2.33,
  2.24,    2.24,    2.24,    2.24,
  2.33,    2.33,    2.33,    2.33,
  2.17,    2.17,    2.17,    2.17,
  2.04,    2.04,    2.04,    2.04,
  2.17,    2.17,    2.17,    2.17,
  2.48,    2.48,    2.48,    2.48,
  2.27,    2.27,    2.27,    2.27,
  2.28,    2.28,    2.28,    2.28,
  2.35,    2.35,    2.35,    2.35,
  2.13,    2.13,    2.13,    2.13,
  2.43,    2.43,    2.43,    2.43,
  2.25,    2.25,    2.25,    2.25,
  2.52,    2.52,    2.52,    2.52,
  2.85,    2.85,    2.85,    2.85,
  2.96,    2.96,    2.96,    2.96,
  2.7,     2.7,     2.7,     2.7,
  2.83,    2.83,    2.83,    2.83,
  3.52,    3.52,    3.52,    3.52,
  3.27,    3.27,    3.27,    3.27,
  3.71,    3.71,    3.71,    3.71,
  3.34,    3.34,    3.34,    3.34,
  3.66,    3.66,    3.66,    3.66,
  2.88,    2.88,    2.88,    2.88,
  3.2,     3.2,     3.2,     3.2,
  3.34,    3.34,    3.34,    3.34,
  4.7,     4.7,     4.7,     4.7,
  4.35,    4.35,    4.35,    4.35,
  3.73,    3.73,    3.73,    3.73,
  4.19,    4.19,    4.19,    4.19,
  3.22,    3.22,    3.22,    3.22,
  3.36,    3.36,    3.36,    3.36,
  3.47,    3.47,    3.47,    3.47,
  2.78,    2.78,    2.78,    2.78,
  3.57,    3.57,    3.57,    3.57,
  2.65,    2.65,    2.65,    2.65,
  2.72,    2.72,    2.72,    2.72,
  2.33,    2.33,    2.33,    2.33,
  1.61,    1.61,    1.61,    1.61,
  2.37,    2.37,    2.37,    2.37,
  2.45,    2.45,    2.45,    2.45,
  1.86,    1.86,    1.86,    1.86,
  1.03,    1.03,    1.03,    1.03,
  1.15,    1.15,    1.15,    1.15,
  1.97,    1.97,    1.97,    1.97,
  2.06,    2.06,    2.06,    2.06,
  2.21,    2.21,    2.21,    2.21,
  2.32,    2.32,    2.32,    2.32,
  2.54,    2.54,    2.54,    2.54,
  2.1,     2.1,     2.1,     2.1,
  2.4,     2.4,     2.4,     2.4,
  2.56,    2.56,    2.56,    2.56,
  2.41,    2.41,    2.41,    2.41,
  2.49,    2.49,    2.49,    2.49,
  2.43,    2.43,    2.43,    2.43,
  2.58,    2.58,    2.58,    2.58,
  2.29,    2.29,    2.29,    2.29,
  2.27,    2.27,    2.27,    2.27,
  2.45,    2.45,    2.45,    2.45,
  2.67,    2.67,    2.67,    2.67,
  2.19,    2.19,    2.19,    2.19,
  2.85,    2.85,    2.85,    2.85,
  2.37,    2.37,    2.37,    2.37,
  2.11,    2.11,    2.11,    2.11,
  2.04,    2.04,    2.04,    2.04,
  2.28,    2.28,    2.28,    2.28,
  2.23,    2.23,    2.23,    2.23,
  2.32,    2.32,    2.32,    2.32,
  2.8,     2.8,     2.8,     2.8,
  2.16,    2.16,    2.16,    2.16,
  2.82,    2.82,    2.82,    2.82,
  3.34,    3.34,    3.34,    3.34,
  3.44,    3.44,    3.44,    3.44,
  4.03,    4.03,    4.03,    4.03,
  3.47,    3.47,    3.47,    3.47,
  3.19,    3.19,    3.19,    3.19,
  3.94,    3.94,    3.94,    3.94,
  1.85,    1.85,    1.85,    1.85,
  2.46,    2.46,    2.46,    2.46,
  2.74,    2.74,    2.74,    2.74,
  2.28,    2.28,    2.28,    2.28,
  3.35,    3.35,    3.35,    3.35,
  3.66,    3.66,    3.66,    3.66,
  3.76,    3.76,    3.76,    3.76,
  4.03,    4.03,    4.03,    4.03,
  2.91,    2.91,    2.91,    2.91,
  2.09,    2.09,    2.09,    2.09,
  1.5,     1.5,     1.5,     1.5,
  0.61,    0.61,    0.61,    0.61,
  1.9,     1.9,     1.9,     1.9,
  2.46,    2.46,    2.46,    2.46,
  2.32,    2.32,    2.32,    2.32,
  1.68,    1.68,    1.68,    1.68,
  1.26,    1.26,    1.26,    1.26,
  1.18,    1.18,    1.18,    1.18,
  1.43,    1.43,    1.43,    1.43,
  1.41,    1.41,    1.41,    1.41,
  1.01,    1.01,    1.01,    1.01,
  1.34,    1.34,    1.34,    1.34,
  1.24,    1.24,    1.24,    1.24,
  1.53,    1.53,    1.53,    1.53,
  2.32,    2.32,    2.32,    2.32,
  2.42,    2.42,    2.42,    2.42,
  3.31,    3.31,    3.31,    3.31,
  3.08,    3.08,    3.08,    3.08,
  3.89,    3.89,    3.89,    3.89,
  4.05,    4.05,    4.05,    4.05,
  3.61,    3.61,    3.61,    3.61,
  3.56,    3.56,    3.56,    3.56,
  3.52,    3.52,    3.52,    3.52,
  3.38,    3.38,    3.38,    3.38,
  3.68,    3.68,    3.68,    3.68,
  3.66,    3.66,    3.66,    3.66,
  3.77,    3.77,    3.77,    3.77,
  4,       4,       4,       4,
  3.58,    3.58,    3.58,    3.58,
  4,       4,       4,       4,
  3.58,    3.58,    3.58,    3.58,
  3.78,    3.78,    3.78,    3.78,
  4.04,    4.04,    4.04,    4.04,
  3.95,    3.95,    3.95,    3.95,
  3.35,    3.35,    3.35,    3.35,
  3.53,    3.53,    3.53,    3.53,
  3.22,    3.22,    3.22,    3.22,
  3.4,     3.4,     3.4,     3.4,
  2.61,    2.61,    2.61,    2.61,
  3.12,    3.12,    3.12,    3.12,
  3.23,    3.23,    3.23,    3.23,
  2.93,    2.93,    2.93,    2.93,
  2.95,    2.95,    2.95,    2.95,
  2.95,    2.95,    2.95,    2.95,
  1.67,    1.67,    1.67,    1.67,
  2,       2,       2,       2,
  2.66,    2.66,    2.66,    2.66,
  2.73,    2.73,    2.73,    2.73,
  2.14,    2.14,    2.14,    2.14,
  2.43,    2.43,    2.43,    2.43,
  1.62,    1.62,    1.62,    1.62,
  1.36,    1.36,    1.36,    1.36,
  1.35,    1.35,    1.35,    1.35,
  1.36,    1.36,    1.36,    1.36,
  1.49,    1.49,    1.49,    1.49,
  1.78,    1.78,    1.78,    1.78,
  1.8,     1.8,     1.8,     1.8,
  2.01,    2.01,    2.01,    2.01,
  1.92,    1.92,    1.92,    1.92,
  1.84,    1.84,    1.84,    1.84,
  1.81,    1.81,    1.81,    1.81,
  1.8,     1.8,     1.8,     1.8,
  1.73,    1.73,    1.73,    1.73,
  2.14,    2.14,    2.14,    2.14,
  1.97,    1.97,    1.97,    1.97,
  1.81,    1.81,    1.81,    1.81,
  1.81,    1.81,    1.81,    1.81,
  2.02,    2.02,    2.02,    2.02,
  1.81,    1.81,    1.81,    1.81,
  1.58,    1.58,    1.58,    1.58,
  1.76,    1.76,    1.76,    1.76,
  1.99,    1.99,    1.99,    1.99,
  1.78,    1.78,    1.78,    1.78,
  2.09,    2.09,    2.09,    2.09,
  1.95,    1.95,    1.95,    1.95,
  2.31,    2.31,    2.31,    2.31,
  2.72,    2.72,    2.72,    2.72,
  2.49,    2.49,    2.49,    2.49,
  3.14,    3.14,    3.14,    3.14,
  2.78,    2.78,    2.78,    2.78,
  2.64,    2.64,    2.64,    2.64,
  2.7,     2.7,     2.7,     2.7,
  2.49,    2.49,    2.49,    2.49,
  3.72,    3.72,    3.72,    3.72,
  3.36,    3.36,    3.36,    3.36,
  4.13,    4.13,    4.13,    4.13,
  3.65,    3.65,    3.65,    3.65,
  3.9,     3.9,     3.9,     3.9,
  4.3,     4.3,     4.3,     4.3,
  3.95,    3.95,    3.95,    3.95,
  3.46,    3.46,    3.46,    3.46,
  3.65,    3.65,    3.65,    3.65,
  3.25,    3.25,    3.25,    3.25,
  3.9,     3.9,     3.9,     3.9,
  0.97,    0.97,    0.97,    0.97,
  0.98,    0.98,    0.98,    0.98,
  0.83,    0.83,    0.83,    0.83,
  0.44,    0.44,    0.44,    0.44,
  0.46,    0.46,    0.46,    0.46,
  0.83,    0.83,    0.83,    0.83,
  0.08,    0.08,    0.08,    0.08,
  1.11,    1.11,    1.11,    1.11,
  0.64,    0.64,    0.64,    0.64,
  1.53,    1.53,    1.53,    1.53,
  1.8,     1.8,     1.8,     1.8,
  1.07,    1.07,    1.07,    1.07,
  1.38,    1.38,    1.38,    1.38,
  1.44,    1.44,    1.44,    1.44,
  1.25,    1.25,    1.25,    1.25,
  1.59,    1.59,    1.59,    1.59,
  1.73,    1.73,    1.73,    1.73,
  2.16,    2.16,    2.16,    2.16,
  2.29,    2.29,    2.29,    2.29,
  1.83,    1.83,    1.83,    1.83,
  1.88,    1.88,    1.88,    1.88,
  1.77,    1.77,    1.77,    1.77,
  1.87,    1.87,    1.87,    1.87,
  2.16,    2.16,    2.16,    2.16,
  1.82,    1.82,    1.82,    1.82,
  2.03,    2.03,    2.03,    2.03,
  2.09,    2.09,    2.09,    2.09,
  2.17,    2.17,    2.17,    2.17,
  2,       2,       2,       2,
  1.83,    1.83,    1.83,    1.83,
  3.05,    3.05,    3.05,    3.05,
  2.53,    2.53,    2.53,    2.53,
  2.61,    2.61,    2.61,    2.61,
  2.39,    2.39,    2.39,    2.39,
  2.7,     2.7,     2.7,     2.7,
  3.32,    3.32,    3.32,    3.32,
  3.54,    3.54,    3.54,    3.54,
  3.63,    3.63,    3.63,    3.63,
  3.62,    3.62,    3.62,    3.62,
  3.2,     3.2,     3.2,     3.2,
  3.39,    3.39,    3.39,    3.39,
  3.84,    3.84,    3.84,    3.84,
  3.25,    3.25,    3.25,    3.25,
  4.08,    4.08,    4.08,    4.08,
  3.73,    3.73,    3.73,    3.73,
  2.81,    2.81,    2.81,    2.81,
  2.75,    2.75,    2.75,    2.75,
  2.85,    2.85,    2.85,    2.85,
  2.03,    2.03,    2.03,    2.03,
  2.42,    2.42,    2.42,    2.42,
  2.64,    2.64,    2.64,    2.64,
  1.55,    1.55,    1.55,    1.55,
  2.14,    2.14,    2.14,    2.14,
  3.11,    3.11,    3.11,    3.11,
  3.36,    3.36,    3.36,    3.36,
  3.19,    3.19,    3.19,    3.19,
  3.46,    3.46,    3.46,    3.46,
  3.24,    3.24,    3.24,    3.24,
  3.29,    3.29,    3.29,    3.29,
  3.1,     3.1,     3.1,     3.1,
  2.85,    2.85,    2.85,    2.85,
  2.35,    2.35,    2.35,    2.35,
  2.6,     2.6,     2.6,     2.6,
  2.25,    2.25,    2.25,    2.25,
  2.49,    2.49,    2.49,    2.49,
  2.28,    2.28,    2.28,    2.28,
  1.94,    1.94,    1.94,    1.94,
  2.05,    2.05,    2.05,    2.05,
  2.01,    2.01,    2.01,    2.01,
  1.96,    1.96,    1.96,    1.96,
  2.08,    2.08,    2.08,    2.08,
  2.19,    2.19,    2.19,    2.19,
  2.32,    2.32,    2.32,    2.32,
  2.33,    2.33,    2.33,    2.33,
  2.79,    2.79,    2.79,    2.79,
  3.16,    3.16,    3.16,    3.16,
  2.95,    2.95,    2.95,    2.95,
  3.12,    3.12,    3.12,    3.12,
  3.71,    3.71,    3.71,    3.71,
  3.75,    3.75,    3.75,    3.75,
  3.84,    3.84,    3.84,    3.84,
  3.94,    3.94,    3.94,    3.94,
  3.51,    3.51,    3.51,    3.51,
  4.74,    4.74,    4.74,    4.74,
  3.69,    3.69,    3.69,    3.69,
  3.42,    3.42,    3.42,    3.42,
  3.71,    3.71,    3.71,    3.71,
  4.41,    4.41,    4.41,    4.41,
  4.28,    4.28,    4.28,    4.28,
  3.6,     3.6,     3.6,     3.6,
  3.56,    3.56,    3.56,    3.56,
  3.3,     3.3,     3.3,     3.3,
  2.81,    2.81,    2.81,    2.81,
  3.82,    3.82,    3.82,    3.82,
  3.36,    3.36,    3.36,    3.36,
  3.11,    3.11,    3.11,    3.11,
  2.65,    2.65,    2.65,    2.65,
  2.6,     2.6,     2.6,     2.6,
  2.13,    2.13,    2.13,    2.13,
  1.98,    1.98,    1.98,    1.98,
  4.1,     4.1,     4.1,     4.1,
  1.36,    1.36,    1.36,    1.36,
  1.09,    1.09,    1.09,    1.09,
  1.58,    1.58,    1.58,    1.58,
  1.86,    1.86,    1.86,    1.86,
  1.83,    1.83,    1.83,    1.83,
  1.94,    1.94,    1.94,    1.94,
  1.88,    1.88,    1.88,    1.88,
  1.88,    1.88,    1.88,    1.88,
  2.23,    2.23,    2.23,    2.23,
  2.34,    2.34,    2.34,    2.34,
  2.17,    2.17,    2.17,    2.17,
  1.93,    1.93,    1.93,    1.93,
  1.71,    1.71,    1.71,    1.71,
  1.92,    1.92,    1.92,    1.92,
  1.93,    1.93,    1.93,    1.93,
  1.64,    1.64,    1.64,    1.64,
  1.78,    1.78,    1.78,    1.78,
  1.8,     1.8,     1.8,     1.8,
  1.96,    1.96,    1.96,    1.96,
  1.95,    1.95,    1.95,    1.95,
  2.12,    2.12,    2.12,    2.12,
  1.78,    1.78,    1.78,    1.78,
  1.58,    1.58,    1.58,    1.58,
  2.05,    2.05,    2.05,    2.05,
  2.01,    2.01,    2.01,    2.01,
  2.58,    2.58,    2.58,    2.58,
  1.55,    1.55,    1.55,    1.55,
  2.23,    2.23,    2.23,    2.23,
  2.46,    2.46,    2.46,    2.46,
  2.49,    2.49,    2.49,    2.49,
  3.18,    3.18,    3.18,    3.18,
  2.97,    2.97,    2.97,    2.97,
  2.8,     2.8,     2.8,     2.8,
  3.14,    3.14,    3.14,    3.14,
  2.94,    2.94,    2.94,    2.94,
  1.94,    1.94,    1.94,    1.94,
  1.37,    1.37,    1.37,    1.37,
  2.63,    2.63,    2.63,    2.63,
  2.8,     2.8,     2.8,     2.8,
  2.2,     2.2,     2.2,     2.2,
  2.42,    2.42,    2.42,    2.42,
  2.01,    2.01,    2.01,    2.01,
  2.14,    2.14,    2.14,    2.14,
  1.91,    1.91,    1.91,    1.91,
  1.54,    1.54,    1.54,    1.54,
  3.39,    3.39,    3.39,    3.39,
  2.85,    2.85,    2.85,    2.85,
  2.6,     2.6,     2.6,     2.6,
  2.37,    2.37,    2.37,    2.37,
  1.6,     1.6,     1.6,     1.6,
  0.94,    0.94,    0.94,    0.94,
  0.79,    0.79,    0.79,    0.79,
  0.54,    0.54,    0.54,    0.54,
  0.59,    0.59,    0.59,    0.59,
  0.78,    0.78,    0.78,    0.78,
  0.5,     0.5,     0.5,     0.5,
  0.66,    0.66,    0.66,    0.66,
  0.77,    0.77,    0.77,    0.77,
  0.84,    0.84,    0.84,    0.84,
  1.07,    1.07,    1.07,    1.07,
  0.86,    0.86,    0.86,    0.86,
  1.11,    1.11,    1.11,    1.11,
  1.13,    1.13,    1.13,    1.13,
  1.27,    1.27,    1.27,    1.27,
  1.58,    1.58,    1.58,    1.58,
  0.22,    0.22,    0.22,    0.22,
  1.06,    1.06,    1.06,    1.06,
  1.67,    1.67,    1.67,    1.67,
  1.32,    1.32,    1.32,    1.32,
  1.08,    1.08,    1.08,    1.08,
  0.68,    0.68,    0.68,    0.68,
  0.58,    0.58,    0.58,    0.58,
  0.57,    0.57,    0.57,    0.57,
  1.21,    1.21,    1.21,    1.21,
  1.36,    1.36,    1.36,    1.36,
  1.4,     1.4,     1.4,     1.4,
  1.56,    1.56,    1.56,    1.56,
  1.15,    1.15,    1.15,    1.15,
  1.84,    1.84,    1.84,    1.84,
  1.17,    1.17,    1.17,    1.17,
  0.82,    0.82,    0.82,    0.82,
  2.36,    2.36,    2.36,    2.36,
  2.48,    2.48,    2.48,    2.48,
  0.18,    0.18,    0.18,    0.18,
  0.72,    0.72,    0.72,    0.72,
  0.24,    0.24,    0.24,    0.24,
  1.45,    1.45,    1.45,    1.45,
  2.13,    2.13,    2.13,    2.13,
  0.91,    0.91,    0.91,    0.91,
  0.66,    0.66,    0.66,    0.66,
  0.81,    0.81,    0.81,    0.81,
  0.7,     0.7,     0.7,     0.7,
  1.06,    1.06,    1.06,    1.06,
  1.76,    1.76,    1.76,    1.76,
  3.16,    3.16,    3.16,    3.16,
  3.24,    3.24,    3.24,    3.24,
  3.24,    3.24,    3.24,    3.24,
  2.81,    2.81,    2.81,    2.81,
  2.47,    2.47,    2.47,    2.47,
  1.79,    1.79,    1.79,    1.79,
  1.96,    1.96,    1.96,    1.96,
  1.37,    1.37,    1.37,    1.37,
  1.43,    1.43,    1.43,    1.43,
  1.32,    1.32,    1.32,    1.32,
  1.97,    1.97,    1.97,    1.97,
  2.22,    2.22,    2.22,    2.22,
  2.14,    2.14,    2.14,    2.14,
  2.09,    2.09,    2.09,    2.09,
  1.92,    1.92,    1.92,    1.92,
  1.67,    1.67,    1.67,    1.67,
  1.83,    1.83,    1.83,    1.83,
  2,       2,       2,       2,
  2.18,    2.18,    2.18,    2.18,
  2.14,    2.14,    2.14,    2.14,
  1.96,    1.96,    1.96,    1.96,
  1.98,    1.98,    1.98,    1.98,
  1.27,    1.27,    1.27,    1.27,
  1.71,    1.71,    1.71,    1.71,
  1.72,    1.72,    1.72,    1.72,
  2.72,    2.72,    2.72,    2.72,
  2.42,    2.42,    2.42,    2.42,
  2.5,     2.5,     2.5,     2.5,
  2.6,     2.6,     2.6,     2.6,
  2.59,    2.59,    2.59,    2.59,
  3.2,     3.2,     3.2,     3.2,
  3.6,     3.6,     3.6,     3.6,
  2.69,    2.69,    2.69,    2.69,
  3.09,    3.09,    3.09,    3.09,
  2.79,    2.79,    2.79,    2.79,
  2.1,     2.1,     2.1,     2.1,
  2.93,    2.93,    2.93,    2.93,
  2.92,    2.92,    2.92,    2.92,
  2.83,    2.83,    2.83,    2.83,
  2.67,    2.67,    2.67,    2.67,
  2.77,    2.77,    2.77,    2.77,
  2.58,    2.58,    2.58,    2.58,
  1.39,    1.39,    1.39,    1.39,
  0.98,    0.98,    0.98,    0.98,
  1.33,    1.33,    1.33,    1.33,
  1.59,    1.59,    1.59,    1.59,
  1.49,    1.49,    1.49,    1.49,
  1.34,    1.34,    1.34,    1.34,
  1.14,    1.14,    1.14,    1.14,
  1.35,    1.35,    1.35,    1.35,
  1.27,    1.27,    1.27,    1.27,
  1.53,    1.53,    1.53,    1.53,
  2.54,    2.54,    2.54,    2.54,
  2.19,    2.19,    2.19,    2.19,
  2.21,    2.21,    2.21,    2.21,
  2.2,     2.2,     2.2,     2.2,
  2.44,    2.44,    2.44,    2.44,
  1.96,    1.96,    1.96,    1.96,
  1.74,    1.74,    1.74,    1.74,
  1.86,    1.86,    1.86,    1.86,
  1.34,    1.34,    1.34,    1.34,
  1.4,     1.4,     1.4,     1.4,
  1.62,    1.62,    1.62,    1.62,
  1.37,    1.37,    1.37,    1.37,
  1.61,    1.61,    1.61,    1.61,
  1.35,    1.35,    1.35,    1.35,
  1.48,    1.48,    1.48,    1.48,
  1.61,    1.61,    1.61,    1.61,
  1.13,    1.13,    1.13,    1.13,
  1.33,    1.33,    1.33,    1.33,
  1.87,    1.87,    1.87,    1.87,
  1.79,    1.79,    1.79,    1.79,
  1.64,    1.64,    1.64,    1.64,
  2.12,    2.12,    2.12,    2.12,
  2.2,     2.2,     2.2,     2.2,
  1.46,    1.46,    1.46,    1.46,
  1.91,    1.91,    1.91,    1.91,
  2.51,    2.51,    2.51,    2.51,
  2.74,    2.74,    2.74,    2.74,
  2.69,    2.69,    2.69,    2.69,
  2.78,    2.78,    2.78,    2.78,
  2.97,    2.97,    2.97,    2.97,
  3.26,    3.26,    3.26,    3.26,
  3.17,    3.17,    3.17,    3.17,
  2.97,    2.97,    2.97,    2.97,
  3.61,    3.61,    3.61,    3.61,
  3.63,    3.63,    3.63,    3.63,
  3.24,    3.24,    3.24,    3.24,
  3.27,    3.27,    3.27,    3.27,
  3.25,    3.25,    3.25,    3.25,
  3.07,    3.07,    3.07,    3.07,
  3.31,    3.31,    3.31,    3.31,
  2.95,    2.95,    2.95,    2.95,
  3.45,    3.45,    3.45,    3.45,
  4.25,    4.25,    4.25,    4.25,
  4.28,    4.28,    4.28,    4.28,
  3.73,    3.73,    3.73,    3.73,
  3.4,     3.4,     3.4,     3.4,
  2.87,    2.87,    2.87,    2.87,
  3.05,    3.05,    3.05,    3.05,
  3.13,    3.13,    3.13,    3.13,
  2.7,     2.7,     2.7,     2.7,
  1.95,    1.95,    1.95,    1.95,
  1.9,     1.9,     1.9,     1.9,
  2.14,    2.14,    2.14,    2.14,
  2.16,    2.16,    2.16,    2.16,
  1.85,    1.85,    1.85,    1.85,
  1.96,    1.96,    1.96,    1.96,
  1.33,    1.33,    1.33,    1.33,
  1.24,    1.24,    1.24,    1.24,
  1.46,    1.46,    1.46,    1.46,
  1.71,    1.71,    1.71,    1.71,
  1.67,    1.67,    1.67,    1.67,
  1.47,    1.47,    1.47,    1.47,
  1.5,     1.5,     1.5,     1.5,
  1.81,    1.81,    1.81,    1.81,
  1.74,    1.74,    1.74,    1.74,
  1.55,    1.55,    1.55,    1.55,
  1.19,    1.19,    1.19,    1.19,
  1.65,    1.65,    1.65,    1.65,
  1.76,    1.76,    1.76,    1.76,
  1.66,    1.66,    1.66,    1.66,
  2.17,    2.17,    2.17,    2.17,
  2.54,    2.54,    2.54,    2.54,
  2.37,    2.37,    2.37,    2.37,
  1.96,    1.96,    1.96,    1.96,
  2.4,     2.4,     2.4,     2.4,
  2.19,    2.19,    2.19,    2.19,
  1.93,    1.93,    1.93,    1.93,
  2.66,    2.66,    2.66,    2.66,
  2.03,    2.03,    2.03,    2.03,
  2.03,    2.03,    2.03,    2.03,
  1.66,    1.66,    1.66,    1.66,
  0.94,    0.94,    0.94,    0.94,
  1.26,    1.26,    1.26,    1.26,
  1.92,    1.92,    1.92,    1.92,
  2.04,    2.04,    2.04,    2.04,
  2.05,    2.05,    2.05,    2.05,
  2.55,    2.55,    2.55,    2.55,
  2.32,    2.32,    2.32,    2.32,
  2.03,    2.03,    2.03,    2.03,
  2.31,    2.31,    2.31,    2.31,
  2.4,     2.4,     2.4,     2.4,
  2.45,    2.45,    2.45,    2.45,
  2.81,    2.81,    2.81,    2.81,
  2.97,    2.97,    2.97,    2.97,
  2.15,    2.15,    2.15,    2.15,
  2,       2,       2,       2,
  1.84,    1.84,    1.84,    1.84,
  2.11,    2.11,    2.11,    2.11,
  2.1,     2.1,     2.1,     2.1,
  2.22,    2.22,    2.22,    2.22,
  2.41,    2.41,    2.41,    2.41,
  2.36,    2.36,    2.36,    2.36,
  1.97,    1.97,    1.97,    1.97,
  1.78,    1.78,    1.78,    1.78,
  1.92,    1.92,    1.92,    1.92,
  1.6,     1.6,     1.6,     1.6,
  1.54,    1.54,    1.54,    1.54,
  1.63,    1.63,    1.63,    1.63,
  1.67,    1.67,    1.67,    1.67,
  1.42,    1.42,    1.42,    1.42,
  1.92,    1.92,    1.92,    1.92,
  2.03,    2.03,    2.03,    2.03,
  2.48,    2.48,    2.48,    2.48,
  1.94,    1.94,    1.94,    1.94,
  2.77,    2.77,    2.77,    2.77,
  1.91,    1.91,    1.91,    1.91,
  1.67,    1.67,    1.67,    1.67,
  1.17,    1.17,    1.17,    1.17,
  2.05,    2.05,    2.05,    2.05,
  1.93,    1.93,    1.93,    1.93,
  1.14,    1.14,    1.14,    1.14,
  1.76,    1.76,    1.76,    1.76,
  1.68,    1.68,    1.68,    1.68,
  2.29,    2.29,    2.29,    2.29,
  2.37,    2.37,    2.37,    2.37,
  2.67,    2.67,    2.67,    2.67,
  3.09,    3.09,    3.09,    3.09,
  2.68,    2.68,    2.68,    2.68,
  1.45,    1.45,    1.45,    1.45,
  1.72,    1.72,    1.72,    1.72,
  1.75,    1.75,    1.75,    1.75,
  1.88,    1.88,    1.88,    1.88,
  1.63,    1.63,    1.63,    1.63,
  2.52,    2.52,    2.52,    2.52,
  2.65,    2.65,    2.65,    2.65,
  2.39,    2.39,    2.39,    2.39,
  2.85,    2.85,    2.85,    2.85,
  2.72,    2.72,    2.72,    2.72,
  2.5,     2.5,     2.5,     2.5,
  2.52,    2.52,    2.52,    2.52,
  2.76,    2.76,    2.76,    2.76,
  2.43,    2.43,    2.43,    2.43,
  2.49,    2.49,    2.49,    2.49,
  2.36,    2.36,    2.36,    2.36,
  2.43,    2.43,    2.43,    2.43,
  2.22,    2.22,    2.22,    2.22,
  2.1,     2.1,     2.1,     2.1,
  2.26,    2.26,    2.26,    2.26,
  2.22,    2.22,    2.22,    2.22,
  2.22,    2.22,    2.22,    2.22,
  2.17,    2.17,    2.17,    2.17,
  2.06,    2.06,    2.06,    2.06,
  2.27,    2.27,    2.27,    2.27,
  1.99,    1.99,    1.99,    1.99,
  1.77,    1.77,    1.77,    1.77,
  1.81,    1.81,    1.81,    1.81,
  1.68,    1.68,    1.68,    1.68,
  1.56,    1.56,    1.56,    1.56,
  1.51,    1.51,    1.51,    1.51,
  1.46,    1.46,    1.46,    1.46,
  1.4,     1.4,     1.4,     1.4,
  1.83,    1.83,    1.83,    1.83,
  2.06,    2.06,    2.06,    2.06,
  2.35,    2.35,    2.35,    2.35,
  2,       2,       2,       2,
  1.52,    1.52,    1.52,    1.52,
  1.74,    1.74,    1.74,    1.74,
  1.78,    1.78,    1.78,    1.78,
  2.1,     2.1,     2.1,     2.1,
  2.06,    2.06,    2.06,    2.06,
  2.83,    2.83,    2.83,    2.83,
  3.55,    3.55,    3.55,    3.55,
  4.03,    4.03,    4.03,    4.03,
  3.71,    3.71,    3.71,    3.71,
  2.64,    2.64,    2.64,    2.64,
  2.95,    2.95,    2.95,    2.95,
  3.21,    3.21,    3.21,    3.21,
  2.84,    2.84,    2.84,    2.84,
  2.95,    2.95,    2.95,    2.95,
  2.71,    2.71,    2.71,    2.71,
  3.21,    3.21,    3.21,    3.21,
  2.83,    2.83,    2.83,    2.83,
  3.54,    3.54,    3.54,    3.54,
  3.67,    3.67,    3.67,    3.67,
  3,       3,       3,       3,
  3.76,    3.76,    3.76,    3.76,
  3.5,     3.5,     3.5,     3.5,
  3.34,    3.34,    3.34,    3.34,
  2.45,    2.45,    2.45,    2.45,
  2.2,     2.2,     2.2,     2.2,
  1.98,    1.98,    1.98,    1.98,
  2.03,    2.03,    2.03,    2.03,
  2.37,    2.37,    2.37,    2.37,
  2.44,    2.44,    2.44,    2.44,
  2.58,    2.58,    2.58,    2.58,
  2.33,    2.33,    2.33,    2.33,
  2.25,    2.25,    2.25,    2.25,
  2.59,    2.59,    2.59,    2.59,
  2.89,    2.89,    2.89,    2.89,
  2.72,    2.72,    2.72,    2.72,
  2.36,    2.36,    2.36,    2.36,
  2.64,    2.64,    2.64,    2.64,
  2.99,    2.99,    2.99,    2.99,
  3.07,    3.07,    3.07,    3.07,
  3.22,    3.22,    3.22,    3.22,
  3.03,    3.03,    3.03,    3.03,
  2.97,    2.97,    2.97,    2.97,
  2.98,    2.98,    2.98,    2.98,
  2.93,    2.93,    2.93,    2.93,
  2.62,    2.62,    2.62,    2.62,
  2.53,    2.53,    2.53,    2.53,
  2.34,    2.34,    2.34,    2.34,
  2.48,    2.48,    2.48,    2.48,
  1.82,    1.82,    1.82,    1.82,
  1.54,    1.54,    1.54,    1.54,
  1.95,    1.95,    1.95,    1.95,
  1.88,    1.88,    1.88,    1.88,
  2.4,     2.4,     2.4,     2.4,
  2.4,     2.4,     2.4,     2.4,
  2.8,     2.8,     2.8,     2.8,
  3.23,    3.23,    3.23,    3.23,
  3.05,    3.05,    3.05,    3.05,
  2.72,    2.72,    2.72,    2.72,
  2.33,    2.33,    2.33,    2.33,
  2.37,    2.37,    2.37,    2.37,
  2.36,    2.36,    2.36,    2.36,
  2.64,    2.64,    2.64,    2.64,
  1.62,    1.62,    1.62,    1.62,
  2.43,    2.43,    2.43,    2.43,
  2.3,     2.3,     2.3,     2.3,
  1.96,    1.96,    1.96,    1.96,
  2.26,    2.26,    2.26,    2.26,
  2.3,     2.3,     2.3,     2.3,
  2.16,    2.16,    2.16,    2.16,
  2.69,    2.69,    2.69,    2.69,
  2.72,    2.72,    2.72,    2.72,
  2.63,    2.63,    2.63,    2.63,
  2.54,    2.54,    2.54,    2.54,
  2.19,    2.19,    2.19,    2.19,
  2.3,     2.3,     2.3,     2.3,
  2.45,    2.45,    2.45,    2.45,
  1.98,    1.98,    1.98,    1.98,
  2.09,    2.09,    2.09,    2.09,
  2.82,    2.82,    2.82,    2.82,
  2.84,    2.84,    2.84,    2.84,
  2.94,    2.94,    2.94,    2.94,
  3.01,    3.01,    3.01,    3.01,
  3.16,    3.16,    3.16,    3.16,
  3.37,    3.37,    3.37,    3.37,
  2.99,    2.99,    2.99,    2.99,
  3.09,    3.09,    3.09,    3.09,
  2.87,    2.87,    2.87,    2.87,
  2.68,    2.68,    2.68,    2.68,
  3.41,    3.41,    3.41,    3.41,
  3.17,    3.17,    3.17,    3.17,
  2.85,    2.85,    2.85,    2.85,
  1.97,    1.97,    1.97,    1.97,
  1.19,    1.19,    1.19,    1.19,
  1.02,    1.02,    1.02,    1.02,
  1.52,    1.52,    1.52,    1.52,
  1.61,    1.61,    1.61,    1.61,
  2.01,    2.01,    2.01,    2.01,
  2.04,    2.04,    2.04,    2.04,
  1.15,    1.15,    1.15,    1.15,
  1.62,    1.62,    1.62,    1.62,
  1.14,    1.14,    1.14,    1.14,
  1.84,    1.84,    1.84,    1.84,
  2.44,    2.44,    2.44,    2.44,
  2.48,    2.48,    2.48,    2.48,
  3.26,    3.26,    3.26,    3.26,
  3.09,    3.09,    3.09,    3.09,
  2.46,    2.46,    2.46,    2.46,
  2.73,    2.73,    2.73,    2.73,
  2.93,    2.93,    2.93,    2.93,
  1.87,    1.87,    1.87,    1.87,
  2.72,    2.72,    2.72,    2.72,
  1.48,    1.48,    1.48,    1.48,
  0.59,    0.59,    0.59,    0.59,
  0.96,    0.96,    0.96,    0.96,
  2.24,    2.24,    2.24,    2.24,
  2.39,    2.39,    2.39,    2.39,
  2.66,    2.66,    2.66,    2.66,
  2.21,    2.21,    2.21,    2.21,
  2.69,    2.69,    2.69,    2.69,
  2.89,    2.89,    2.89,    2.89,
  2.11,    2.11,    2.11,    2.11,
  2.17,    2.17,    2.17,    2.17,
  1.85,    1.85,    1.85,    1.85,
  1.64,    1.64,    1.64,    1.64,
  1.36,    1.36,    1.36,    1.36,
  1.16,    1.16,    1.16,    1.16,
  1.11,    1.11,    1.11,    1.11,
  1.44,    1.44,    1.44,    1.44,
  1.25,    1.25,    1.25,    1.25,
  1.51,    1.51,    1.51,    1.51,
  1.49,    1.49,    1.49,    1.49,
  1.43,    1.43,    1.43,    1.43,
  1.72,    1.72,    1.72,    1.72,
  1.82,    1.82,    1.82,    1.82,
  1.95,    1.95,    1.95,    1.95,
  1.31,    1.31,    1.31,    1.31,
  1.02,    1.02,    1.02,    1.02,
  1.16,    1.16,    1.16,    1.16,
  1.25,    1.25,    1.25,    1.25,
  0.94,    0.94,    0.94,    0.94,
  0.61,    0.61,    0.61,    0.61,
  0.33,    0.33,    0.33,    0.33,
  0.27,    0.27,    0.27,    0.27,
  0.18,    0.18,    0.18,    0.18,
  0.67,    0.67,    0.67,    0.67,
  0.57,    0.57,    0.57,    0.57,
  0.38,    0.38,    0.38,    0.38,
  0.76,    0.76,    0.76,    0.76,
  0.29,    0.29,    0.29,    0.29,
  0.98,    0.98,    0.98,    0.98,
  1.48,    1.48,    1.48,    1.48,
  1.21,    1.21,    1.21,    1.21,
  1.64,    1.64,    1.64,    1.64,
  1.87,    1.87,    1.87,    1.87,
  1.38,    1.38,    1.38,    1.38,
  1.34,    1.34,    1.34,    1.34,
  1.53,    1.53,    1.53,    1.53,
  1.59,    1.59,    1.59,    1.59,
  1.94,    1.94,    1.94,    1.94,
  2.75,    2.75,    2.75,    2.75,
  1.98,    1.98,    1.98,    1.98,
  2.6,     2.6,     2.6,     2.6,
  2.25,    2.25,    2.25,    2.25,
  1.26,    1.26,    1.26,    1.26,
  1.96,    1.96,    1.96,    1.96,
  2.37,    2.37,    2.37,    2.37,
  1.43,    1.43,    1.43,    1.43,
  2.08,    2.08,    2.08,    2.08,
  1.46,    1.46,    1.46,    1.46,
  0.86,    0.86,    0.86,    0.86,
  1.96,    1.96,    1.96,    1.96,
  1.5,     1.5,     1.5,     1.5,
  1.04,    1.04,    1.04,    1.04,
  0.81,    0.81,    0.81,    0.81,
  1.35,    1.35,    1.35,    1.35,
  1.19,    1.19,    1.19,    1.19,
  0.8,     0.8,     0.8,     0.8,
  1.15,    1.15,    1.15,    1.15,
  1.34,    1.34,    1.34,    1.34,
  1.5,     1.5,     1.5,     1.5,
  0.89,    0.89,    0.89,    0.89,
  0.41,    0.41,    0.41,    0.41,
  1.13,    1.13,    1.13,    1.13,
  1.22,    1.22,    1.22,    1.22,
  1.78,    1.78,    1.78,    1.78,
  1.91,    1.91,    1.91,    1.91,
  1.76,    1.76,    1.76,    1.76,
  1.72,    1.72,    1.72,    1.72,
  1.78,    1.78,    1.78,    1.78,
  1.33,    1.33,    1.33,    1.33,
  1.38,    1.38,    1.38,    1.38,
  0.42,    0.42,    0.42,    0.42,
  0.94,    0.94,    0.94,    0.94,
  1.39,    1.39,    1.39,    1.39,
  1.38,    1.38,    1.38,    1.38,
  1.2,     1.2,     1.2,     1.2,
  1.37,    1.37,    1.37,    1.37,
  2.82,    2.82,    2.82,    2.82,
  2.9,     2.9,     2.9,     2.9,
  2.88,    2.88,    2.88,    2.88,
  3.73,    3.73,    3.73,    3.73,
  2.82,    2.82,    2.82,    2.82,
  3.18,    3.18,    3.18,    3.18,
  3.06,    3.06,    3.06,    3.06,
  3.01,    3.01,    3.01,    3.01,
  3.03,    3.03,    3.03,    3.03,
  2.42,    2.42,    2.42,    2.42,
  2.41,    2.41,    2.41,    2.41,
  2.62,    2.62,    2.62,    2.62,
  2.54,    2.54,    2.54,    2.54,
  2.67,    2.67,    2.67,    2.67,
  3.35,    3.35,    3.35,    3.35,
  2.68,    2.68,    2.68,    2.68,
  2.79,    2.79,    2.79,    2.79,
  3.5,     3.5,     3.5,     3.5,
  2.99,    2.99,    2.99,    2.99,
  3.17,    3.17,    3.17,    3.17,
  2.17,    2.17,    2.17,    2.17,
  2.05,    2.05,    2.05,    2.05,
  2.14,    2.14,    2.14,    2.14,
  2.14,    2.14,    2.14,    2.14,
  1.86,    1.86,    1.86,    1.86,
  2.35,    2.35,    2.35,    2.35,
  2.19,    2.19,    2.19,    2.19,
  2.16,    2.16,    2.16,    2.16,
  1.1,     1.1,     1.1,     1.1,
  0.63,    0.63,    0.63,    0.63,
  1.25,    1.25,    1.25,    1.25,
  1.66,    1.66,    1.66,    1.66,
  1.85,    1.85,    1.85,    1.85,
  1.73,    1.73,    1.73,    1.73,
  1.64,    1.64,    1.64,    1.64,
  1.71,    1.71,    1.71,    1.71,
  1.55,    1.55,    1.55,    1.55,
  1.13,    1.13,    1.13,    1.13,
  1.34,    1.34,    1.34,    1.34,
  1.26,    1.26,    1.26,    1.26,
  1.54,    1.54,    1.54,    1.54,
  0.89,    0.89,    0.89,    0.89,
  0.54,    0.54,    0.54,    0.54,
  0.78,    0.78,    0.78,    0.78,
  1.15,    1.15,    1.15,    1.15,
  1.44,    1.44,    1.44,    1.44,
  1.32,    1.32,    1.32,    1.32,
  1.08,    1.08,    1.08,    1.08,
  1.69,    1.69,    1.69,    1.69,
  1.76,    1.76,    1.76,    1.76,
  2.23,    2.23,    2.23,    2.23,
  2,       2,       2,       2,
  3.14,    3.14,    3.14,    3.14,
  2.68,    2.68,    2.68,    2.68,
  1.18,    1.18,    1.18,    1.18,
  1.43,    1.43,    1.43,    1.43,
  2.65,    2.65,    2.65,    2.65,
  2.95,    2.95,    2.95,    2.95,
  2.94,    2.94,    2.94,    2.94,
  2.12,    2.12,    2.12,    2.12,
  1.9,     1.9,     1.9,     1.9,
  2.91,    2.91,    2.91,    2.91,
  1.97,    1.97,    1.97,    1.97,
  1.8,     1.8,     1.8,     1.8,
  1.01,    1.01,    1.01,    1.01,
  1.05,    1.05,    1.05,    1.05,
  0.93,    0.93,    0.93,    0.93,
  1.64,    1.64,    1.64,    1.64,
  1.01,    1.01,    1.01,    1.01,
  0.52,    0.52,    0.52,    0.52,
  0.37,    0.37,    0.37,    0.37,
  1.05,    1.05,    1.05,    1.05,
  1.33,    1.33,    1.33,    1.33,
  1.81,    1.81,    1.81,    1.81,
  1.99,    1.99,    1.99,    1.99,
  2.12,    2.12,    2.12,    2.12,
  2.17,    2.17,    2.17,    2.17,
  2.06,    2.06,    2.06,    2.06,
  1.79,    1.79,    1.79,    1.79,
  1.73,    1.73,    1.73,    1.73,
  1.82,    1.82,    1.82,    1.82,
  1.92,    1.92,    1.92,    1.92,
  2.01,    2.01,    2.01,    2.01,
  2.13,    2.13,    2.13,    2.13,
  2.3,     2.3,     2.3,     2.3,
  2.42,    2.42,    2.42,    2.42,
  1.69,    1.69,    1.69,    1.69,
  1.57,    1.57,    1.57,    1.57,
  1.68,    1.68,    1.68,    1.68,
  1.5,     1.5,     1.5,     1.5,
  1.76,    1.76,    1.76,    1.76,
  1.91,    1.91,    1.91,    1.91,
  2.14,    2.14,    2.14,    2.14,
  2.48,    2.48,    2.48,    2.48,
  2.4,     2.4,     2.4,     2.4,
  2.4,     2.4,     2.4,     2.4,
  2.57,    2.57,    2.57,    2.57,
  2.32,    2.32,    2.32,    2.32,
  2.07,    2.07,    2.07,    2.07,
  2.8,     2.8,     2.8,     2.8,
  2.54,    2.54,    2.54,    2.54,
  2.54,    2.54,    2.54,    2.54,
  3.02,    3.02,    3.02,    3.02,
  3.29,    3.29,    3.29,    3.29,
  3.51,    3.51,    3.51,    3.51,
  3.31,    3.31,    3.31,    3.31,
  3.66,    3.66,    3.66,    3.66,
  4.13,    4.13,    4.13,    4.13,
  3.81,    3.81,    3.81,    3.81,
  3.05,    3.05,    3.05,    3.05,
  3.31,    3.31,    3.31,    3.31,
  3.22,    3.22,    3.22,    3.22,
  3.38,    3.38,    3.38,    3.38,
  2.46,    2.46,    2.46,    2.46,
  3.54,    3.54,    3.54,    3.54,
  2.18,    2.18,    2.18,    2.18,
  2.43,    2.43,    2.43,    2.43,
  2.49,    2.49,    2.49,    2.49,
  1.88,    1.88,    1.88,    1.88,
  1.43,    1.43,    1.43,    1.43,
  1.41,    1.41,    1.41,    1.41,
  0.98,    0.98,    0.98,    0.98,
  1.54,    1.54,    1.54,    1.54,
  1.36,    1.36,    1.36,    1.36,
  1.48,    1.48,    1.48,    1.48,
  1.46,    1.46,    1.46,    1.46,
  1.4,     1.4,     1.4,     1.4,
  1.5,     1.5,     1.5,     1.5,
  1.17,    1.17,    1.17,    1.17,
  1.45,    1.45,    1.45,    1.45,
  1.4,     1.4,     1.4,     1.4,
  1.38,    1.38,    1.38,    1.38,
  1.54,    1.54,    1.54,    1.54,
  1.48,    1.48,    1.48,    1.48,
  1.18,    1.18,    1.18,    1.18,
  1.28,    1.28,    1.28,    1.28,
  1.1,     1.1,     1.1,     1.1,
  1.26,    1.26,    1.26,    1.26,
  1.87,    1.87,    1.87,    1.87,
  1.97,    1.97,    1.97,    1.97,
  2.3,     2.3,     2.3,     2.3,
  2.24,    2.24,    2.24,    2.24,
  2.53,    2.53,    2.53,    2.53,
  2.36,    2.36,    2.36,    2.36,
  3.16,    3.16,    3.16,    3.16,
  2.88,    2.88,    2.88,    2.88,
  3.33,    3.33,    3.33,    3.33,
  2.92,    2.92,    2.92,    2.92,
  2.96,    2.96,    2.96,    2.96,
  2.88,    2.88,    2.88,    2.88,
  3.48,    3.48,    3.48,    3.48,
  3.09,    3.09,    3.09,    3.09,
  2.7,     2.7,     2.7,     2.7,
  3.73,    3.73,    3.73,    3.73,
  3.69,    3.69,    3.69,    3.69,
  3.52,    3.52,    3.52,    3.52,
  3.4,     3.4,     3.4,     3.4,
  3.18,    3.18,    3.18,    3.18,
  2.68,    2.68,    2.68,    2.68,
  2.45,    2.45,    2.45,    2.45,
  2.48,    2.48,    2.48,    2.48,
  2.14,    2.14,    2.14,    2.14,
  1.56,    1.56,    1.56,    1.56,
  1.09,    1.09,    1.09,    1.09,
  1.66,    1.66,    1.66,    1.66,
  1.73,    1.73,    1.73,    1.73,
  1.92,    1.92,    1.92,    1.92,
  1.81,    1.81,    1.81,    1.81,
  1.84,    1.84,    1.84,    1.84,
  1.34,    1.34,    1.34,    1.34,
  1.1,     1.1,     1.1,     1.1,
  0.91,    0.91,    0.91,    0.91,
  0.08,    0.08,    0.08,    0.08,
  0.53,    0.53,    0.53,    0.53,
  0.6,     0.6,     0.6,     0.6,
  0.68,    0.68,    0.68,    0.68,
  1.24,    1.24,    1.24,    1.24,
  1.32,    1.32,    1.32,    1.32,
  1.2,     1.2,     1.2,     1.2,
  1.09,    1.09,    1.09,    1.09,
  1.01,    1.01,    1.01,    1.01,
  0.76,    0.76,    0.76,    0.76,
  0.74,    0.74,    0.74,    0.74,
  0.92,    0.92,    0.92,    0.92,
  0.72,    0.72,    0.72,    0.72,
  0.75,    0.75,    0.75,    0.75,
  0.67,    0.67,    0.67,    0.67,
  0.9,     0.9,     0.9,     0.9,
  0.77,    0.77,    0.77,    0.77,
  1.78,    1.78,    1.78,    1.78,
  1.6,     1.6,     1.6,     1.6,
  1.38,    1.38,    1.38,    1.38,
  1.71,    1.71,    1.71,    1.71,
  2.08,    2.08,    2.08,    2.08,
  0.96,    0.96,    0.96,    0.96,
  1.38,    1.38,    1.38,    1.38,
  1.2,     1.2,     1.2,     1.2,
  1.96,    1.96,    1.96,    1.96,
  1.86,    1.86,    1.86,    1.86,
  2.42,    2.42,    2.42,    2.42,
  1.77,    1.77,    1.77,    1.77,
  1.95,    1.95,    1.95,    1.95,
  2.21,    2.21,    2.21,    2.21,
  2.52,    2.52,    2.52,    2.52,
  2.19,    2.19,    2.19,    2.19,
  1.68,    1.68,    1.68,    1.68,
  1.84,    1.84,    1.84,    1.84,
  2.13,    2.13,    2.13,    2.13,
  1.51,    1.51,    1.51,    1.51,
  0.94,    0.94,    0.94,    0.94,
  2.34,    2.34,    2.34,    2.34,
  1.97,    1.97,    1.97,    1.97,
  2.19,    2.19,    2.19,    2.19,
  2,       2,       2,       2,
  2.2,     2.2,     2.2,     2.2,
  2.21,    2.21,    2.21,    2.21,
  2.39,    2.39,    2.39,    2.39,
  2.75,    2.75,    2.75,    2.75,
  2.43,    2.43,    2.43,    2.43,
  2.23,    2.23,    2.23,    2.23,
  2.5,     2.5,     2.5,     2.5,
  2.79,    2.79,    2.79,    2.79,
  2.53,    2.53,    2.53,    2.53,
  2.62,    2.62,    2.62,    2.62,
  2.45,    2.45,    2.45,    2.45,
  2.61,    2.61,    2.61,    2.61,
  2.44,    2.44,    2.44,    2.44,
  2.33,    2.33,    2.33,    2.33,
  2.38,    2.38,    2.38,    2.38,
  2.45,    2.45,    2.45,    2.45,
  2.34,    2.34,    2.34,    2.34,
  2.17,    2.17,    2.17,    2.17,
  2.05,    2.05,    2.05,    2.05,
  2.08,    2.08,    2.08,    2.08,
  2.36,    2.36,    2.36,    2.36,
  2.34,    2.34,    2.34,    2.34,
  3.2,     3.2,     3.2,     3.2,
  3.04,    3.04,    3.04,    3.04,
  2.28,    2.28,    2.28,    2.28,
  2.66,    2.66,    2.66,    2.66,
  3.06,    3.06,    3.06,    3.06,
  3.31,    3.31,    3.31,    3.31,
  3.89,    3.89,    3.89,    3.89,
  3.34,    3.34,    3.34,    3.34,
  3.42,    3.42,    3.42,    3.42,
  3.55,    3.55,    3.55,    3.55,
  3.23,    3.23,    3.23,    3.23,
  3.56,    3.56,    3.56,    3.56,
  2.62,    2.62,    2.62,    2.62,
  2.23,    2.23,    2.23,    2.23,
  1.83,    1.83,    1.83,    1.83,
  3.03,    3.03,    3.03,    3.03,
  3.41,    3.41,    3.41,    3.41,
  4.23,    4.23,    4.23,    4.23,
  4.2,     4.2,     4.2,     4.2,
  4,       4,       4,       4,
  3.13,    3.13,    3.13,    3.13,
  3.34,    3.34,    3.34,    3.34,
  3.45,    3.45,    3.45,    3.45,
  2.47,    2.47,    2.47,    2.47,
  2.2,     2.2,     2.2,     2.2,
  1.83,    1.83,    1.83,    1.83,
  2.12,    2.12,    2.12,    2.12,
  1.97,    1.97,    1.97,    1.97,
  2.19,    2.19,    2.19,    2.19,
  2.26,    2.26,    2.26,    2.26,
  2.26,    2.26,    2.26,    2.26,
  1.93,    1.93,    1.93,    1.93,
  2.03,    2.03,    2.03,    2.03,
  2.15,    2.15,    2.15,    2.15,
  1.84,    1.84,    1.84,    1.84,
  1.91,    1.91,    1.91,    1.91,
  2.12,    2.12,    2.12,    2.12,
  2,       2,       2,       2,
  1.82,    1.82,    1.82,    1.82,
  1.84,    1.84,    1.84,    1.84,
  1.97,    1.97,    1.97,    1.97,
  1.78,    1.78,    1.78,    1.78,
  1.25,    1.25,    1.25,    1.25,
  1.57,    1.57,    1.57,    1.57,
  1.69,    1.69,    1.69,    1.69,
  1.48,    1.48,    1.48,    1.48,
  1.58,    1.58,    1.58,    1.58,
  1.53,    1.53,    1.53,    1.53,
  1.61,    1.61,    1.61,    1.61,
  1.78,    1.78,    1.78,    1.78,
  1.69,    1.69,    1.69,    1.69,
  1.49,    1.49,    1.49,    1.49,
  2.5,     2.5,     2.5,     2.5,
  3.14,    3.14,    3.14,    3.14,
  2.88,    2.88,    2.88,    2.88,
  3.58,    3.58,    3.58,    3.58,
  3.48,    3.48,    3.48,    3.48,
  3.08,    3.08,    3.08,    3.08,
  2.95,    2.95,    2.95,    2.95,
  2.84,    2.84,    2.84,    2.84,
  2.62,    2.62,    2.62,    2.62,
  2.77,    2.77,    2.77,    2.77,
  2.94,    2.94,    2.94,    2.94,
  1.52,    1.52,    1.52,    1.52,
  0.39,    0.39,    0.39,    0.39,
  0.84,    0.84,    0.84,    0.84,
  1.26,    1.26,    1.26,    1.26,
  1.23,    1.23,    1.23,    1.23,
  1.05,    1.05,    1.05,    1.05,
  2.07,    2.07,    2.07,    2.07,
  2.77,    2.77,    2.77,    2.77,
  3.02,    3.02,    3.02,    3.02,
  2.73,    2.73,    2.73,    2.73,
  2.77,    2.77,    2.77,    2.77,
  2.42,    2.42,    2.42,    2.42,
  2.73,    2.73,    2.73,    2.73,
  2.6,     2.6,     2.6,     2.6,
  2.42,    2.42,    2.42,    2.42,
  2.44,    2.44,    2.44,    2.44,
  2.27,    2.27,    2.27,    2.27,
  2.47,    2.47,    2.47,    2.47,
  2.28,    2.28,    2.28,    2.28,
  2.09,    2.09,    2.09,    2.09,
  2.47,    2.47,    2.47,    2.47,
  2.32,    2.32,    2.32,    2.32,
  2.18,    2.18,    2.18,    2.18,
  2.03,    2.03,    2.03,    2.03,
  2,       2,       2,       2,
  2.3,     2.3,     2.3,     2.3,
  2.34,    2.34,    2.34,    2.34,
  2.44,    2.44,    2.44,    2.44,
  2.47,    2.47,    2.47,    2.47,
  2.35,    2.35,    2.35,    2.35,
  2.25,    2.25,    2.25,    2.25,
  2.17,    2.17,    2.17,    2.17,
  2.14,    2.14,    2.14,    2.14,
  2.32,    2.32,    2.32,    2.32,
  2.75,    2.75,    2.75,    2.75,
  2.84,    2.84,    2.84,    2.84,
  2.69,    2.69,    2.69,    2.69,
  2.45,    2.45,    2.45,    2.45,
  2.83,    2.83,    2.83,    2.83,
  3.44,    3.44,    3.44,    3.44,
  3.72,    3.72,    3.72,    3.72,
  3.44,    3.44,    3.44,    3.44,
  2.95,    2.95,    2.95,    2.95,
  2.18,    2.18,    2.18,    2.18,
  2.92,    2.92,    2.92,    2.92,
  2.25,    2.25,    2.25,    2.25,
  2.16,    2.16,    2.16,    2.16,
  3.39,    3.39,    3.39,    3.39,
  2.41,    2.41,    2.41,    2.41,
  1.46,    1.46,    1.46,    1.46,
  2.98,    2.98,    2.98,    2.98,
  2.31,    2.31,    2.31,    2.31,
  1.96,    1.96,    1.96,    1.96,
  2.02,    2.02,    2.02,    2.02,
  2.32,    2.32,    2.32,    2.32,
  2.31,    2.31,    2.31,    2.31,
  2.3,     2.3,     2.3,     2.3,
  1.96,    1.96,    1.96,    1.96,
  1.85,    1.85,    1.85,    1.85,
  2.14,    2.14,    2.14,    2.14,
  1.95,    1.95,    1.95,    1.95,
  2.76,    2.76,    2.76,    2.76,
  3.57,    3.57,    3.57,    3.57,
  2.89,    2.89,    2.89,    2.89,
  2.38,    2.38,    2.38,    2.38,
  1.66,    1.66,    1.66,    1.66,
  1.77,    1.77,    1.77,    1.77,
  1.94,    1.94,    1.94,    1.94,
  1.63,    1.63,    1.63,    1.63,
  1.73,    1.73,    1.73,    1.73,
  1.38,    1.38,    1.38,    1.38,
  1.53,    1.53,    1.53,    1.53,
  1.71,    1.71,    1.71,    1.71,
  1.47,    1.47,    1.47,    1.47,
  1.53,    1.53,    1.53,    1.53,
  1.86,    1.86,    1.86,    1.86,
  1.46,    1.46,    1.46,    1.46,
  1.52,    1.52,    1.52,    1.52,
  1.46,    1.46,    1.46,    1.46,
  1.61,    1.61,    1.61,    1.61,
  1.85,    1.85,    1.85,    1.85,
  1.74,    1.74,    1.74,    1.74,
  1.82,    1.82,    1.82,    1.82,
  1.32,    1.32,    1.32,    1.32,
  1.54,    1.54,    1.54,    1.54,
  1.57,    1.57,    1.57,    1.57,
  2,       2,       2,       2,
  2.23,    2.23,    2.23,    2.23,
  1.95,    1.95,    1.95,    1.95,
  1.79,    1.79,    1.79,    1.79,
  2.63,    2.63,    2.63,    2.63,
  2.58,    2.58,    2.58,    2.58,
  2.2,     2.2,     2.2,     2.2,
  0.3,     0.3,     0.3,     0.3,
  1.76,    1.76,    1.76,    1.76,
  1.56,    1.56,    1.56,    1.56,
  2.01,    2.01,    2.01,    2.01,
  1.71,    1.71,    1.71,    1.71,
  1.67,    1.67,    1.67,    1.67,
  1.51,    1.51,    1.51,    1.51,
  2.77,    2.77,    2.77,    2.77,
  2.87,    2.87,    2.87,    2.87,
  2.16,    2.16,    2.16,    2.16,
  2.1,     2.1,     2.1,     2.1,
  1.87,    1.87,    1.87,    1.87,
  1.65,    1.65,    1.65,    1.65,
  1.53,    1.53,    1.53,    1.53,
  1.65,    1.65,    1.65,    1.65,
  1.71,    1.71,    1.71,    1.71,
  2.09,    2.09,    2.09,    2.09,
  1.75,    1.75,    1.75,    1.75,
  1.87,    1.87,    1.87,    1.87,
  2.21,    2.21,    2.21,    2.21,
  1.56,    1.56,    1.56,    1.56,
  1.47,    1.47,    1.47,    1.47,
  1.02,    1.02,    1.02,    1.02,
  1.36,    1.36,    1.36,    1.36,
  1.63,    1.63,    1.63,    1.63,
  1.67,    1.67,    1.67,    1.67,
  1.17,    1.17,    1.17,    1.17,
  1.36,    1.36,    1.36,    1.36,
  1.44,    1.44,    1.44,    1.44,
  1.34,    1.34,    1.34,    1.34,
  1.41,    1.41,    1.41,    1.41,
  1.49,    1.49,    1.49,    1.49,
  1.67,    1.67,    1.67,    1.67,
  1.37,    1.37,    1.37,    1.37,
  1.31,    1.31,    1.31,    1.31,
  1.35,    1.35,    1.35,    1.35,
  1.73,    1.73,    1.73,    1.73,
  2.24,    2.24,    2.24,    2.24,
  2.42,    2.42,    2.42,    2.42,
  2.52,    2.52,    2.52,    2.52,
  2.28,    2.28,    2.28,    2.28,
  2.04,    2.04,    2.04,    2.04,
  2.17,    2.17,    2.17,    2.17,
  1.79,    1.79,    1.79,    1.79,
  2.58,    2.58,    2.58,    2.58,
  2.61,    2.61,    2.61,    2.61,
  2.64,    2.64,    2.64,    2.64,
  3.23,    3.23,    3.23,    3.23,
  3.13,    3.13,    3.13,    3.13,
  3.74,    3.74,    3.74,    3.74,
  3.71,    3.71,    3.71,    3.71,
  2.65,    2.65,    2.65,    2.65,
  2.69,    2.69,    2.69,    2.69,
  3.01,    3.01,    3.01,    3.01,
  2.78,    2.78,    2.78,    2.78,
  2.6,     2.6,     2.6,     2.6,
  2.91,    2.91,    2.91,    2.91,
  2.12,    2.12,    2.12,    2.12,
  2.02,    2.02,    2.02,    2.02,
  1.32,    1.32,    1.32,    1.32,
  1.26,    1.26,    1.26,    1.26,
  1.84,    1.84,    1.84,    1.84,
  1.63,    1.63,    1.63,    1.63,
  1.67,    1.67,    1.67,    1.67,
  1.74,    1.74,    1.74,    1.74,
  1.72,    1.72,    1.72,    1.72,
  1.72,    1.72,    1.72,    1.72,
  2.16,    2.16,    2.16,    2.16,
  2.11,    2.11,    2.11,    2.11,
  2.13,    2.13,    2.13,    2.13,
  2.24,    2.24,    2.24,    2.24,
  2.65,    2.65,    2.65,    2.65,
  2.52,    2.52,    2.52,    2.52,
  2.64,    2.64,    2.64,    2.64,
  2.64,    2.64,    2.64,    2.64,
  2.5,     2.5,     2.5,     2.5,
  2.37,    2.37,    2.37,    2.37,
  2.1,     2.1,     2.1,     2.1,
  1.93,    1.93,    1.93,    1.93,
  1.94,    1.94,    1.94,    1.94,
  1.7,     1.7,     1.7,     1.7,
  1.67,    1.67,    1.67,    1.67,
  1.82,    1.82,    1.82,    1.82,
  1.44,    1.44,    1.44,    1.44,
  1.7,     1.7,     1.7,     1.7,
  1.34,    1.34,    1.34,    1.34,
  1.8,     1.8,     1.8,     1.8,
  1.5,     1.5,     1.5,     1.5,
  1.8,     1.8,     1.8,     1.8,
  1.64,    1.64,    1.64,    1.64,
  1.66,    1.66,    1.66,    1.66,
  1.87,    1.87,    1.87,    1.87,
  2.7,     2.7,     2.7,     2.7,
  2.77,    2.77,    2.77,    2.77,
  2.97,    2.97,    2.97,    2.97,
  3.49,    3.49,    3.49,    3.49,
  2.11,    2.11,    2.11,    2.11,
  1.55,    1.55,    1.55,    1.55,
  1.15,    1.15,    1.15,    1.15,
  1.39,    1.39,    1.39,    1.39,
  1.42,    1.42,    1.42,    1.42,
  1.97,    1.97,    1.97,    1.97,
  2.76,    2.76,    2.76,    2.76,
  3.02,    3.02,    3.02,    3.02,
  3.07,    3.07,    3.07,    3.07,
  1.56,    1.56,    1.56,    1.56,
  1.28,    1.28,    1.28,    1.28,
  0.74,    0.74,    0.74,    0.74,
  1.16,    1.16,    1.16,    1.16,
  1.3,     1.3,     1.3,     1.3,
  1.44,    1.44,    1.44,    1.44,
  1.58,    1.58,    1.58,    1.58,
  1.64,    1.64,    1.64,    1.64,
  1.62,    1.62,    1.62,    1.62,
  1.33,    1.33,    1.33,    1.33,
  2.05,    2.05,    2.05,    2.05,
  1.84,    1.84,    1.84,    1.84,
  1.96,    1.96,    1.96,    1.96,
  1.76,    1.76,    1.76,    1.76,
  1.86,    1.86,    1.86,    1.86,
  1.75,    1.75,    1.75,    1.75,
  1.66,    1.66,    1.66,    1.66,
  1.61,    1.61,    1.61,    1.61,
  1.69,    1.69,    1.69,    1.69,
  1.61,    1.61,    1.61,    1.61,
  1.72,    1.72,    1.72,    1.72,
  1.99,    1.99,    1.99,    1.99,
  2.64,    2.64,    2.64,    2.64,
  1.89,    1.89,    1.89,    1.89,
  1.55,    1.55,    1.55,    1.55,
  1.87,    1.87,    1.87,    1.87,
  2.12,    2.12,    2.12,    2.12,
  2.19,    2.19,    2.19,    2.19,
  2,       2,       2,       2,
  2.84,    2.84,    2.84,    2.84,
  2.47,    2.47,    2.47,    2.47,
  2.8,     2.8,     2.8,     2.8,
  2.31,    2.31,    2.31,    2.31,
  2.45,    2.45,    2.45,    2.45,
  4.83,    4.83,    4.83,    4.83,
  3.31,    3.31,    3.31,    3.31,
  3.4,     3.4,     3.4,     3.4,
  4.03,    4.03,    4.03,    4.03,
  4.36,    4.36,    4.36,    4.36,
  3.45,    3.45,    3.45,    3.45,
  4.02,    4.02,    4.02,    4.02,
  5.21,    5.21,    5.21,    5.21,
  5.29,    5.29,    5.29,    5.29,
  6.25,    6.25,    6.25,    6.25,
  6.08,    6.08,    6.08,    6.08,
  5.45,    5.45,    5.45,    5.45,
  5.47,    5.47,    5.47,    5.47,
  6.12,    6.12,    6.12,    6.12,
  5.72,    5.72,    5.72,    5.72,
  5.21,    5.21,    5.21,    5.21,
  4.81,    4.81,    4.81,    4.81,
  4.31,    4.31,    4.31,    4.31,
  3.46,    3.46,    3.46,    3.46,
  3.45,    3.45,    3.45,    3.45,
  3.2,     3.2,     3.2,     3.2,
  2.69,    2.69,    2.69,    2.69,
  2.45,    2.45,    2.45,    2.45,
  2.37,    2.37,    2.37,    2.37,
  2.27,    2.27,    2.27,    2.27,
  2.39,    2.39,    2.39,    2.39,
  2.13,    2.13,    2.13,    2.13,
  1.93,    1.93,    1.93,    1.93,
  2.08,    2.08,    2.08,    2.08,
  1.99,    1.99,    1.99,    1.99,
  2.18,    2.18,    2.18,    2.18,
  2.64,    2.64,    2.64,    2.64,
  2.22,    2.22,    2.22,    2.22,
  2.59,    2.59,    2.59,    2.59,
  2.87,    2.87,    2.87,    2.87,
  3.12,    3.12,    3.12,    3.12,
  2.87,    2.87,    2.87,    2.87,
  3.12,    3.12,    3.12,    3.12,
  3.5,     3.5,     3.5,     3.5,
  3.2,     3.2,     3.2,     3.2,
  4.16,    4.16,    4.16,    4.16,
  4.02,    4.02,    4.02,    4.02,
  4.12,    4.12,    4.12,    4.12,
  3.92,    3.92,    3.92,    3.92,
  3.81,    3.81,    3.81,    3.81,
  3.36,    3.36,    3.36,    3.36,
  4.2,     4.2,     4.2,     4.2,
  3.48,    3.48,    3.48,    3.48,
  4.01,    4.01,    4.01,    4.01,
  4.03,    4.03,    4.03,    4.03,
  4.2,     4.2,     4.2,     4.2,
  4.06,    4.06,    4.06,    4.06,
  3.99,    3.99,    3.99,    3.99,
  3.04,    3.04,    3.04,    3.04,
  3.55,    3.55,    3.55,    3.55,
  3.03,    3.03,    3.03,    3.03,
  2.93,    2.93,    2.93,    2.93,
  3.56,    3.56,    3.56,    3.56,
  3.67,    3.67,    3.67,    3.67,
  3.34,    3.34,    3.34,    3.34,
  2.99,    2.99,    2.99,    2.99,
  1.94,    1.94,    1.94,    1.94,
  1.65,    1.65,    1.65,    1.65,
  1.86,    1.86,    1.86,    1.86,
  2.31,    2.31,    2.31,    2.31,
  1.63,    1.63,    1.63,    1.63,
  1.97,    1.97,    1.97,    1.97,
  2.18,    2.18,    2.18,    2.18,
  2.59,    2.59,    2.59,    2.59,
  2.91,    2.91,    2.91,    2.91,
  3.62,    3.62,    3.62,    3.62,
  2.71,    2.71,    2.71,    2.71,
  2.99,    2.99,    2.99,    2.99,
  3.55,    3.55,    3.55,    3.55,
  3.4,     3.4,     3.4,     3.4,
  3.62,    3.62,    3.62,    3.62,
  3.76,    3.76,    3.76,    3.76,
  3.84,    3.84,    3.84,    3.84,
  4.52,    4.52,    4.52,    4.52,
  3.84,    3.84,    3.84,    3.84,
  5.16,    5.16,    5.16,    5.16,
  4.44,    4.44,    4.44,    4.44,
  4.19,    4.19,    4.19,    4.19,
  3.71,    3.71,    3.71,    3.71,
  3.68,    3.68,    3.68,    3.68,
  3.87,    3.87,    3.87,    3.87,
  3.79,    3.79,    3.79,    3.79,
  3.67,    3.67,    3.67,    3.67,
  3.56,    3.56,    3.56,    3.56,
  4.29,    4.29,    4.29,    4.29,
  4.62,    4.62,    4.62,    4.62,
  4.34,    4.34,    4.34,    4.34,
  4.67,    4.67,    4.67,    4.67,
  5.23,    5.23,    5.23,    5.23,
  5.91,    5.91,    5.91,    5.91,
  5.25,    5.25,    5.25,    5.25,
  4.25,    4.25,    4.25,    4.25,
  5.45,    5.45,    5.45,    5.45,
  5.26,    5.26,    5.26,    5.26,
  4.24,    4.24,    4.24,    4.24,
  4.61,    4.61,    4.61,    4.61,
  4.55,    4.55,    4.55,    4.55,
  5.28,    5.28,    5.28,    5.28,
  4.5,     4.5,     4.5,     4.5,
  5.46,    5.46,    5.46,    5.46,
  5.78,    5.78,    5.78,    5.78,
  4.94,    4.94,    4.94,    4.94,
  4.55,    4.55,    4.55,    4.55,
  4.53,    4.53,    4.53,    4.53,
  4.51,    4.51,    4.51,    4.51,
  3.74,    3.74,    3.74,    3.74,
  4.2,     4.2,     4.2,     4.2,
  3.31,    3.31,    3.31,    3.31,
  3.09,    3.09,    3.09,    3.09,
  2.3,     2.3,     2.3,     2.3,
  2.13,    2.13,    2.13,    2.13,
  2.19,    2.19,    2.19,    2.19,
  1.99,    1.99,    1.99,    1.99,
  2.02,    2.02,    2.02,    2.02,
  2.09,    2.09,    2.09,    2.09,
  1.84,    1.84,    1.84,    1.84,
  1.92,    1.92,    1.92,    1.92,
  1.94,    1.94,    1.94,    1.94,
  1.89,    1.89,    1.89,    1.89,
  1.88,    1.88,    1.88,    1.88,
  1.68,    1.68,    1.68,    1.68,
  2.04,    2.04,    2.04,    2.04,
  2.12,    2.12,    2.12,    2.12,
  2.2,     2.2,     2.2,     2.2,
  2.04,    2.04,    2.04,    2.04,
  2.01,    2.01,    2.01,    2.01,
  1.89,    1.89,    1.89,    1.89,
  1.9,     1.9,     1.9,     1.9,
  1.74,    1.74,    1.74,    1.74,
  1.51,    1.51,    1.51,    1.51,
  1.52,    1.52,    1.52,    1.52,
  1.54,    1.54,    1.54,    1.54,
  1.78,    1.78,    1.78,    1.78,
  1.84,    1.84,    1.84,    1.84,
  3.13,    3.13,    3.13,    3.13,
  3.04,    3.04,    3.04,    3.04,
  3.01,    3.01,    3.01,    3.01,
  3.35,    3.35,    3.35,    3.35,
  3.3,     3.3,     3.3,     3.3,
  2.7,     2.7,     2.7,     2.7,
  3.1,     3.1,     3.1,     3.1,
  3.25,    3.25,    3.25,    3.25,
  3.61,    3.61,    3.61,    3.61,
  4.05,    4.05,    4.05,    4.05,
  4.27,    4.27,    4.27,    4.27,
  3.75,    3.75,    3.75,    3.75,
  4.4,     4.4,     4.4,     4.4,
  3.27,    3.27,    3.27,    3.27,
  2.87,    2.87,    2.87,    2.87,
  3.18,    3.18,    3.18,    3.18,
  2.69,    2.69,    2.69,    2.69,
  3.42,    3.42,    3.42,    3.42,
  4.08,    4.08,    4.08,    4.08,
  4.06,    4.06,    4.06,    4.06,
  2.58,    2.58,    2.58,    2.58,
  2.6,     2.6,     2.6,     2.6,
  1.9,     1.9,     1.9,     1.9,
  2.06,    2.06,    2.06,    2.06,
  2,       2,       2,       2,
  1.51,    1.51,    1.51,    1.51,
  2.09,    2.09,    2.09,    2.09,
  2.02,    2.02,    2.02,    2.02,
  1.12,    1.12,    1.12,    1.12,
  0.77,    0.77,    0.77,    0.77,
  0.93,    0.93,    0.93,    0.93,
  0.68,    0.68,    0.68,    0.68,
  0.82,    0.82,    0.82,    0.82,
  1.93,    1.93,    1.93,    1.93,
  1.87,    1.87,    1.87,    1.87,
  1.47,    1.47,    1.47,    1.47,
  1.41,    1.41,    1.41,    1.41,
  1.71,    1.71,    1.71,    1.71,
  1.06,    1.06,    1.06,    1.06,
  1.72,    1.72,    1.72,    1.72,
  2.16,    2.16,    2.16,    2.16,
  1.79,    1.79,    1.79,    1.79,
  1.29,    1.29,    1.29,    1.29,
  1.4,     1.4,     1.4,     1.4,
  0.43,    0.43,    0.43,    0.43,
  1.12,    1.12,    1.12,    1.12,
  1.33,    1.33,    1.33,    1.33,
  1.7,     1.7,     1.7,     1.7,
  2.03,    2.03,    2.03,    2.03,
  2.24,    2.24,    2.24,    2.24,
  1.51,    1.51,    1.51,    1.51,
  1.14,    1.14,    1.14,    1.14,
  1.01,    1.01,    1.01,    1.01,
  1.82,    1.82,    1.82,    1.82,
  1.82,    1.82,    1.82,    1.82,
  1.71,    1.71,    1.71,    1.71,
  1.96,    1.96,    1.96,    1.96,
  1.79,    1.79,    1.79,    1.79,
  1.74,    1.74,    1.74,    1.74,
  1.98,    1.98,    1.98,    1.98,
  2.3,     2.3,     2.3,     2.3,
  1.78,    1.78,    1.78,    1.78,
  1.77,    1.77,    1.77,    1.77,
  1.55,    1.55,    1.55,    1.55,
  1.66,    1.66,    1.66,    1.66,
  2.1,     2.1,     2.1,     2.1,
  1.65,    1.65,    1.65,    1.65,
  1.61,    1.61,    1.61,    1.61,
  0.94,    0.94,    0.94,    0.94,
  0.64,    0.64,    0.64,    0.64,
  0.39,    0.39,    0.39,    0.39,
  0.26,    0.26,    0.26,    0.26,
  1.61,    1.61,    1.61,    1.61,
  1.8,     1.8,     1.8,     1.8,
  1.64,    1.64,    1.64,    1.64,
  2.2,     2.2,     2.2,     2.2,
  2.47,    2.47,    2.47,    2.47,
  2.52,    2.52,    2.52,    2.52,
  2.45,    2.45,    2.45,    2.45,
  2.65,    2.65,    2.65,    2.65,
  2.44,    2.44,    2.44,    2.44,
  2.63,    2.63,    2.63,    2.63,
  2.58,    2.58,    2.58,    2.58,
  2.41,    2.41,    2.41,    2.41,
  2.48,    2.48,    2.48,    2.48,
  2.7,     2.7,     2.7,     2.7,
  2.45,    2.45,    2.45,    2.45,
  2.59,    2.59,    2.59,    2.59,
  2.57,    2.57,    2.57,    2.57,
  2.65,    2.65,    2.65,    2.65,
  2.62,    2.62,    2.62,    2.62,
  2.64,    2.64,    2.64,    2.64,
  2.41,    2.41,    2.41,    2.41,
  2.46,    2.46,    2.46,    2.46,
  2.48,    2.48,    2.48,    2.48,
  2.25,    2.25,    2.25,    2.25,
  2.17,    2.17,    2.17,    2.17,
  2.08,    2.08,    2.08,    2.08,
  1.99,    1.99,    1.99,    1.99,
  1.67,    1.67,    1.67,    1.67,
  2.24,    2.24,    2.24,    2.24,
  1.83,    1.83,    1.83,    1.83,
  2.66,    2.66,    2.66,    2.66,
  2.46,    2.46,    2.46,    2.46,
  2.34,    2.34,    2.34,    2.34,
  2.24,    2.24,    2.24,    2.24,
  1.59,    1.59,    1.59,    1.59,
  1.63,    1.63,    1.63,    1.63,
  1.74,    1.74,    1.74,    1.74,
  1.84,    1.84,    1.84,    1.84,
  1.51,    1.51,    1.51,    1.51,
  2.02,    2.02,    2.02,    2.02,
  2.92,    2.92,    2.92,    2.92,
  3.51,    3.51,    3.51,    3.51,
  4.1,     4.1,     4.1,     4.1,
  3.83,    3.83,    3.83,    3.83,
  3.88,    3.88,    3.88,    3.88,
  3.25,    3.25,    3.25,    3.25,
  3.69,    3.69,    3.69,    3.69,
  3.19,    3.19,    3.19,    3.19,
  2.3,     2.3,     2.3,     2.3,
  2.14,    2.14,    2.14,    2.14,
  1.73,    1.73,    1.73,    1.73,
  2.1,     2.1,     2.1,     2.1,
  0.51,    0.51,    0.51,    0.51,
  1.12,    1.12,    1.12,    1.12,
  1.49,    1.49,    1.49,    1.49,
  1.95,    1.95,    1.95,    1.95,
  1.75,    1.75,    1.75,    1.75,
  1.99,    1.99,    1.99,    1.99,
  1.65,    1.65,    1.65,    1.65,
  1.61,    1.61,    1.61,    1.61,
  1.74,    1.74,    1.74,    1.74,
  1.75,    1.75,    1.75,    1.75,
  1.86,    1.86,    1.86,    1.86,
  2.06,    2.06,    2.06,    2.06,
  2.03,    2.03,    2.03,    2.03,
  1.96,    1.96,    1.96,    1.96,
  2.07,    2.07,    2.07,    2.07,
  2.33,    2.33,    2.33,    2.33,
  2.84,    2.84,    2.84,    2.84,
  2.8,     2.8,     2.8,     2.8,
  3.28,    3.28,    3.28,    3.28,
  3.44,    3.44,    3.44,    3.44,
  4.25,    4.25,    4.25,    4.25,
  3.17,    3.17,    3.17,    3.17,
  2.52,    2.52,    2.52,    2.52,
  2.82,    2.82,    2.82,    2.82,
  3.83,    3.83,    3.83,    3.83,
  4.31,    4.31,    4.31,    4.31,
  5,       5,       5,       5,
  4.6,     4.6,     4.6,     4.6,
  5.05,    5.05,    5.05,    5.05,
  5.15,    5.15,    5.15,    5.15,
  5.23,    5.23,    5.23,    5.23,
  5.57,    5.57,    5.57,    5.57,
  5.35,    5.35,    5.35,    5.35,
  2.7,     2.7,     2.7,     2.7,
  3,       3,       3,       3,
  3.28,    3.28,    3.28,    3.28,
  3.57,    3.57,    3.57,    3.57,
  4.02,    4.02,    4.02,    4.02,
  3.8,     3.8,     3.8,     3.8,
  3.9,     3.9,     3.9,     3.9,
  3.95,    3.95,    3.95,    3.95,
  3.55,    3.55,    3.55,    3.55,
  3.1,     3.1,     3.1,     3.1,
  2.82,    2.82,    2.82,    2.82,
  2.39,    2.39,    2.39,    2.39,
  1.99,    1.99,    1.99,    1.99,
  2.47,    2.47,    2.47,    2.47,
  2.23,    2.23,    2.23,    2.23,
  1.56,    1.56,    1.56,    1.56,
  1.62,    1.62,    1.62,    1.62,
  2.05,    2.05,    2.05,    2.05,
  1.8,     1.8,     1.8,     1.8,
  1.78,    1.78,    1.78,    1.78,
  1.73,    1.73,    1.73,    1.73,
  2.18,    2.18,    2.18,    2.18,
  2.42,    2.42,    2.42,    2.42,
  2.14,    2.14,    2.14,    2.14,
  1.58,    1.58,    1.58,    1.58,
  1.63,    1.63,    1.63,    1.63,
  1.7,     1.7,     1.7,     1.7,
  1.63,    1.63,    1.63,    1.63,
  1.71,    1.71,    1.71,    1.71,
  1.8,     1.8,     1.8,     1.8,
  1.33,    1.33,    1.33,    1.33,
  0.79,    0.79,    0.79,    0.79,
  1.61,    1.61,    1.61,    1.61,
  1.44,    1.44,    1.44,    1.44,
  1.59,    1.59,    1.59,    1.59,
  1.66,    1.66,    1.66,    1.66,
  1.58,    1.58,    1.58,    1.58,
  1.63,    1.63,    1.63,    1.63,
  1.24,    1.24,    1.24,    1.24,
  1.61,    1.61,    1.61,    1.61,
  2.37,    2.37,    2.37,    2.37,
  1.99,    1.99,    1.99,    1.99,
  1.97,    1.97,    1.97,    1.97,
  2.41,    2.41,    2.41,    2.41,
  2.49,    2.49,    2.49,    2.49,
  2.31,    2.31,    2.31,    2.31,
  1.67,    1.67,    1.67,    1.67,
  2.11,    2.11,    2.11,    2.11,
  2.47,    2.47,    2.47,    2.47,
  2.75,    2.75,    2.75,    2.75,
  2.73,    2.73,    2.73,    2.73,
  2.29,    2.29,    2.29,    2.29,
  2.25,    2.25,    2.25,    2.25,
  2.39,    2.39,    2.39,    2.39,
  2.3,     2.3,     2.3,     2.3,
  2.01,    2.01,    2.01,    2.01,
  1.9,     1.9,     1.9,     1.9,
  2.22,    2.22,    2.22,    2.22,
  2.11,    2.11,    2.11,    2.11,
  2.12,    2.12,    2.12,    2.12,
  1.77,    1.77,    1.77,    1.77,
  1.38,    1.38,    1.38,    1.38,
  1.37,    1.37,    1.37,    1.37,
  1.46,    1.46,    1.46,    1.46,
  1.42,    1.42,    1.42,    1.42,
  1.54,    1.54,    1.54,    1.54,
  1.47,    1.47,    1.47,    1.47,
  1.71,    1.71,    1.71,    1.71,
  1.74,    1.74,    1.74,    1.74,
  1.66,    1.66,    1.66,    1.66,
  1.78,    1.78,    1.78,    1.78,
  1.79,    1.79,    1.79,    1.79,
  1.92,    1.92,    1.92,    1.92,
  1.33,    1.33,    1.33,    1.33,
  0.9,     0.9,     0.9,     0.9,
  1.37,    1.37,    1.37,    1.37,
  1.82,    1.82,    1.82,    1.82,
  1.76,    1.76,    1.76,    1.76,
  1.45,    1.45,    1.45,    1.45,
  1.38,    1.38,    1.38,    1.38,
  1.61,    1.61,    1.61,    1.61,
  1.53,    1.53,    1.53,    1.53,
  1.35,    1.35,    1.35,    1.35,
  2.38,    2.38,    2.38,    2.38,
  2.04,    2.04,    2.04,    2.04,
  1.6,     1.6,     1.6,     1.6,
  1.71,    1.71,    1.71,    1.71,
  2.11,    2.11,    2.11,    2.11,
  2.21,    2.21,    2.21,    2.21,
  2.44,    2.44,    2.44,    2.44,
  2.6,     2.6,     2.6,     2.6,
  2.59,    2.59,    2.59,    2.59,
  2.94,    2.94,    2.94,    2.94,
  3.31,    3.31,    3.31,    3.31,
  3.19,    3.19,    3.19,    3.19,
  2.92,    2.92,    2.92,    2.92,
  2.86,    2.86,    2.86,    2.86,
  2.86,    2.86,    2.86,    2.86,
  2.14,    2.14,    2.14,    2.14,
  2.2,     2.2,     2.2,     2.2,
  2.29,    2.29,    2.29,    2.29,
  1.88,    1.88,    1.88,    1.88,
  1.98,    1.98,    1.98,    1.98,
  1.85,    1.85,    1.85,    1.85,
  1.39,    1.39,    1.39,    1.39,
  0.95,    0.95,    0.95,    0.95,
  1,       1,       1,       1,
  1.57,    1.57,    1.57,    1.57,
  1.01,    1.01,    1.01,    1.01,
  1.73,    1.73,    1.73,    1.73,
  1.48,    1.48,    1.48,    1.48,
  1.54,    1.54,    1.54,    1.54,
  1.98,    1.98,    1.98,    1.98,
  1.9,     1.9,     1.9,     1.9,
  1.81,    1.81,    1.81,    1.81,
  2.27,    2.27,    2.27,    2.27,
  1.82,    1.82,    1.82,    1.82,
  1.57,    1.57,    1.57,    1.57,
  1.34,    1.34,    1.34,    1.34,
  1.65,    1.65,    1.65,    1.65,
  1.89,    1.89,    1.89,    1.89,
  2.04,    2.04,    2.04,    2.04,
  2.02,    2.02,    2.02,    2.02,
  1.52,    1.52,    1.52,    1.52,
  1.44,    1.44,    1.44,    1.44,
  1.93,    1.93,    1.93,    1.93,
  1.86,    1.86,    1.86,    1.86,
  2.27,    2.27,    2.27,    2.27,
  2.53,    2.53,    2.53,    2.53,
  2.67,    2.67,    2.67,    2.67,
  2.98,    2.98,    2.98,    2.98,
  3.54,    3.54,    3.54,    3.54,
  3.37,    3.37,    3.37,    3.37,
  3.16,    3.16,    3.16,    3.16,
  2.64,    2.64,    2.64,    2.64,
  2.37,    2.37,    2.37,    2.37,
  2.31,    2.31,    2.31,    2.31,
  1.51,    1.51,    1.51,    1.51,
  2.48,    2.48,    2.48,    2.48,
  2.19,    2.19,    2.19,    2.19,
  2.11,    2.11,    2.11,    2.11,
  2.15,    2.15,    2.15,    2.15,
  2.39,    2.39,    2.39,    2.39,
  1.67,    1.67,    1.67,    1.67,
  2.21,    2.21,    2.21,    2.21,
  2.02,    2.02,    2.02,    2.02,
  1.73,    1.73,    1.73,    1.73,
  1.82,    1.82,    1.82,    1.82,
  1.35,    1.35,    1.35,    1.35,
  1.35,    1.35,    1.35,    1.35,
  1.12,    1.12,    1.12,    1.12,
  1.34,    1.34,    1.34,    1.34,
  1.33,    1.33,    1.33,    1.33,
  1.53,    1.53,    1.53,    1.53,
  1.75,    1.75,    1.75,    1.75,
  1.67,    1.67,    1.67,    1.67,
  2.21,    2.21,    2.21,    2.21,
  1.91,    1.91,    1.91,    1.91,
  2.07,    2.07,    2.07,    2.07,
  2.51,    2.51,    2.51,    2.51,
  2.63,    2.63,    2.63,    2.63,
  2.35,    2.35,    2.35,    2.35,
  2.24,    2.24,    2.24,    2.24,
  2.63,    2.63,    2.63,    2.63,
  2.77,    2.77,    2.77,    2.77,
  2.77,    2.77,    2.77,    2.77,
  2.88,    2.88,    2.88,    2.88,
  3.07,    3.07,    3.07,    3.07,
  2.78,    2.78,    2.78,    2.78,
  2.46,    2.46,    2.46,    2.46,
  2.52,    2.52,    2.52,    2.52,
  2.81,    2.81,    2.81,    2.81,
  2.33,    2.33,    2.33,    2.33,
  2.2,     2.2,     2.2,     2.2,
  2.26,    2.26,    2.26,    2.26,
  2.04,    2.04,    2.04,    2.04,
  3,       3,       3,       3,
  3.15,    3.15,    3.15,    3.15,
  3.49,    3.49,    3.49,    3.49,
  4.28,    4.28,    4.28,    4.28,
  3.39,    3.39,    3.39,    3.39,
  3.3,     3.3,     3.3,     3.3,
  3.69,    3.69,    3.69,    3.69,
  3.74,    3.74,    3.74,    3.74,
  3.5,     3.5,     3.5,     3.5,
  3.49,    3.49,    3.49,    3.49,
  3.89,    3.89,    3.89,    3.89,
  3.14,    3.14,    3.14,    3.14,
  2.89,    2.89,    2.89,    2.89,
  2.78,    2.78,    2.78,    2.78,
  3.15,    3.15,    3.15,    3.15,
  2.68,    2.68,    2.68,    2.68,
  2.82,    2.82,    2.82,    2.82,
  2.8,     2.8,     2.8,     2.8,
  2.86,    2.86,    2.86,    2.86,
  3.23,    3.23,    3.23,    3.23,
  2.93,    2.93,    2.93,    2.93,
  3.06,    3.06,    3.06,    3.06,
  3.29,    3.29,    3.29,    3.29,
  2.5,     2.5,     2.5,     2.5,
  2.18,    2.18,    2.18,    2.18,
  1.96,    1.96,    1.96,    1.96,
  2.59,    2.59,    2.59,    2.59,
  3.16,    3.16,    3.16,    3.16,
  3.04,    3.04,    3.04,    3.04,
  2.76,    2.76,    2.76,    2.76,
  2.72,    2.72,    2.72,    2.72,
  2.92,    2.92,    2.92,    2.92,
  3.05,    3.05,    3.05,    3.05,
  3.37,    3.37,    3.37,    3.37,
  2.82,    2.82,    2.82,    2.82,
  2.78,    2.78,    2.78,    2.78,
  2.59,    2.59,    2.59,    2.59,
  2.26,    2.26,    2.26,    2.26,
  2,       2,       2,       2,
  1.91,    1.91,    1.91,    1.91,
  2.16,    2.16,    2.16,    2.16,
  1.29,    1.29,    1.29,    1.29,
  1.11,    1.11,    1.11,    1.11,
  2.01,    2.01,    2.01,    2.01,
  1.37,    1.37,    1.37,    1.37,
  0.18,    0.18,    0.18,    0.18,
  0.81,    0.81,    0.81,    0.81,
  1.73,    1.73,    1.73,    1.73,
  1.58,    1.58,    1.58,    1.58,
  2.52,    2.52,    2.52,    2.52,
  3.2,     3.2,     3.2,     3.2,
  3.16,    3.16,    3.16,    3.16,
  4.23,    4.23,    4.23,    4.23,
  3.71,    3.71,    3.71,    3.71,
  2.89,    2.89,    2.89,    2.89,
  3.48,    3.48,    3.48,    3.48,
  3.26,    3.26,    3.26,    3.26,
  3.74,    3.74,    3.74,    3.74,
  3.74,    3.74,    3.74,    3.74,
  3.96,    3.96,    3.96,    3.96,
  3.66,    3.66,    3.66,    3.66,
  3.83,    3.83,    3.83,    3.83,
  3.54,    3.54,    3.54,    3.54,
  3.35,    3.35,    3.35,    3.35,
  4.05,    4.05,    4.05,    4.05,
  3.93,    3.93,    3.93,    3.93,
  2.42,    2.42,    2.42,    2.42,
  3.11,    3.11,    3.11,    3.11,
  3.92,    3.92,    3.92,    3.92,
  3.03,    3.03,    3.03,    3.03,
  3.52,    3.52,    3.52,    3.52,
  3.65,    3.65,    3.65,    3.65,
  3.08,    3.08,    3.08,    3.08,
  2.5,     2.5,     2.5,     2.5,
  2.04,    2.04,    2.04,    2.04,
  1.95,    1.95,    1.95,    1.95,
  2.34,    2.34,    2.34,    2.34,
  2.74,    2.74,    2.74,    2.74,
  2.98,    2.98,    2.98,    2.98,
  3.11,    3.11,    3.11,    3.11,
  3.32,    3.32,    3.32,    3.32,
  3.52,    3.52,    3.52,    3.52,
  3.63,    3.63,    3.63,    3.63,
  3.68,    3.68,    3.68,    3.68,
  3.22,    3.22,    3.22,    3.22,
  3.07,    3.07,    3.07,    3.07,
  3.19,    3.19,    3.19,    3.19,
  3.22,    3.22,    3.22,    3.22,
  3.2,     3.2,     3.2,     3.2,
  3.33,    3.33,    3.33,    3.33,
  3.63,    3.63,    3.63,    3.63,
  3.55,    3.55,    3.55,    3.55,
  3.18,    3.18,    3.18,    3.18,
  3.08,    3.08,    3.08,    3.08,
  2.93,    2.93,    2.93,    2.93,
  2.93,    2.93,    2.93,    2.93,
  2.61,    2.61,    2.61,    2.61,
  2.8,     2.8,     2.8,     2.8,
  3.1,     3.1,     3.1,     3.1,
  2.97,    2.97,    2.97,    2.97,
  3.2,     3.2,     3.2,     3.2,
  2.81,    2.81,    2.81,    2.81,
  3.71,    3.71,    3.71,    3.71,
  4.23,    4.23,    4.23,    4.23,
  4.61,    4.61,    4.61,    4.61,
  5.27,    5.27,    5.27,    5.27,
  5.04,    5.04,    5.04,    5.04,
  4.89,    4.89,    4.89,    4.89,
  4.92,    4.92,    4.92,    4.92,
  4.62,    4.62,    4.62,    4.62,
  4.6,     4.6,     4.6,     4.6,
  4.4,     4.4,     4.4,     4.4,
  4.19,    4.19,    4.19,    4.19,
  5.03,    5.03,    5.03,    5.03,
  4.56,    4.56,    4.56,    4.56,
  4.54,    4.54,    4.54,    4.54,
  4.6,     4.6,     4.6,     4.6,
  4.4,     4.4,     4.4,     4.4,
  4.76,    4.76,    4.76,    4.76,
  3.7,     3.7,     3.7,     3.7,
  3.49,    3.49,    3.49,    3.49,
  3.42,    3.42,    3.42,    3.42,
  2.65,    2.65,    2.65,    2.65,
  2.7,     2.7,     2.7,     2.7,
  2.61,    2.61,    2.61,    2.61,
  2.9,     2.9,     2.9,     2.9,
  3.13,    3.13,    3.13,    3.13,
  3.43,    3.43,    3.43,    3.43,
  3.35,    3.35,    3.35,    3.35,
  3.21,    3.21,    3.21,    3.21,
  2.94,    2.94,    2.94,    2.94,
  2.86,    2.86,    2.86,    2.86,
  3.18,    3.18,    3.18,    3.18,
  3.23,    3.23,    3.23,    3.23,
  3.14,    3.14,    3.14,    3.14,
  2.67,    2.67,    2.67,    2.67,
  2.88,    2.88,    2.88,    2.88,
  2.9,     2.9,     2.9,     2.9,
  2.98,    2.98,    2.98,    2.98,
  2.8,     2.8,     2.8,     2.8,
  2.89,    2.89,    2.89,    2.89,
  2.64,    2.64,    2.64,    2.64,
  2.62,    2.62,    2.62,    2.62,
  2.5,     2.5,     2.5,     2.5,
  3.14,    3.14,    3.14,    3.14,
  3.7,     3.7,     3.7,     3.7,
  3.52,    3.52,    3.52,    3.52,
  2.83,    2.83,    2.83,    2.83,
  3.26,    3.26,    3.26,    3.26,
  3.83,    3.83,    3.83,    3.83,
  4.42,    4.42,    4.42,    4.42,
  4.52,    4.52,    4.52,    4.52,
  4.62,    4.62,    4.62,    4.62,
  5.25,    5.25,    5.25,    5.25,
  4.44,    4.44,    4.44,    4.44,
  4.49,    4.49,    4.49,    4.49,
  4.34,    4.34,    4.34,    4.34,
  5.11,    5.11,    5.11,    5.11,
  4.54,    4.54,    4.54,    4.54,
  4.97,    4.97,    4.97,    4.97,
  4.82,    4.82,    4.82,    4.82,
  4.26,    4.26,    4.26,    4.26,
  4.1,     4.1,     4.1,     4.1,
  4.29,    4.29,    4.29,    4.29,
  3.98,    3.98,    3.98,    3.98,
  4.31,    4.31,    4.31,    4.31,
  3.81,    3.81,    3.81,    3.81,
  4.38,    4.38,    4.38,    4.38,
  3.43,    3.43,    3.43,    3.43,
  3.09,    3.09,    3.09,    3.09,
  2.74,    2.74,    2.74,    2.74,
  2.6,     2.6,     2.6,     2.6,
  2.63,    2.63,    2.63,    2.63,
  2.61,    2.61,    2.61,    2.61,
  2.65,    2.65,    2.65,    2.65,
  2.86,    2.86,    2.86,    2.86,
  2.9,     2.9,     2.9,     2.9,
  3,       3,       3,       3,
  3.01,    3.01,    3.01,    3.01,
  3.01,    3.01,    3.01,    3.01,
  3.04,    3.04,    3.04,    3.04,
  2.73,    2.73,    2.73,    2.73,
  2.78,    2.78,    2.78,    2.78,
  2.69,    2.69,    2.69,    2.69,
  2.3,     2.3,     2.3,     2.3,
  2.6,     2.6,     2.6,     2.6,
  2.72,    2.72,    2.72,    2.72,
  2.98,    2.98,    2.98,    2.98,
  2.51,    2.51,    2.51,    2.51,
  2.97,    2.97,    2.97,    2.97,
  2.73,    2.73,    2.73,    2.73,
  3.04,    3.04,    3.04,    3.04,
  3.32,    3.32,    3.32,    3.32,
  2.87,    2.87,    2.87,    2.87,
  2.91,    2.91,    2.91,    2.91,
  3.09,    3.09,    3.09,    3.09,
  2.6,     2.6,     2.6,     2.6,
  2.82,    2.82,    2.82,    2.82,
  2.64,    2.64,    2.64,    2.64,
  3.48,    3.48,    3.48,    3.48,
  3.22,    3.22,    3.22,    3.22,
  3.11,    3.11,    3.11,    3.11,
  3.52,    3.52,    3.52,    3.52,
  3.28,    3.28,    3.28,    3.28,
  3.03,    3.03,    3.03,    3.03,
  2.83,    2.83,    2.83,    2.83,
  2.29,    2.29,    2.29,    2.29,
  2.96,    2.96,    2.96,    2.96,
  2.55,    2.55,    2.55,    2.55,
  2.71,    2.71,    2.71,    2.71,
  2.44,    2.44,    2.44,    2.44,
  1.93,    1.93,    1.93,    1.93,
  2.27,    2.27,    2.27,    2.27,
  1.96,    1.96,    1.96,    1.96,
  2.35,    2.35,    2.35,    2.35,
  2.11,    2.11,    2.11,    2.11,
  1.75,    1.75,    1.75,    1.75,
  1.92,    1.92,    1.92,    1.92,
  2.27,    2.27,    2.27,    2.27,
  2.66,    2.66,    2.66,    2.66,
  2.71,    2.71,    2.71,    2.71,
  2.79,    2.79,    2.79,    2.79,
  2.84,    2.84,    2.84,    2.84,
  2.35,    2.35,    2.35,    2.35,
  2.48,    2.48,    2.48,    2.48,
  2.52,    2.52,    2.52,    2.52,
  2.6,     2.6,     2.6,     2.6,
  2.72,    2.72,    2.72,    2.72,
  2.81,    2.81,    2.81,    2.81,
  2.64,    2.64,    2.64,    2.64,
  2.27,    2.27,    2.27,    2.27,
  2.49,    2.49,    2.49,    2.49,
  2.52,    2.52,    2.52,    2.52,
  2.95,    2.95,    2.95,    2.95,
  2.95,    2.95,    2.95,    2.95,
  2.85,    2.85,    2.85,    2.85,
  2.4,     2.4,     2.4,     2.4,
  2.63,    2.63,    2.63,    2.63,
  2.31,    2.31,    2.31,    2.31,
  1.36,    1.36,    1.36,    1.36,
  1.07,    1.07,    1.07,    1.07,
  1.05,    1.05,    1.05,    1.05,
  1.07,    1.07,    1.07,    1.07,
  1.13,    1.13,    1.13,    1.13,
  1.53,    1.53,    1.53,    1.53,
  1.12,    1.12,    1.12,    1.12,
  1.25,    1.25,    1.25,    1.25,
  1.85,    1.85,    1.85,    1.85,
  1,       1,       1,       1,
  0.99,    0.99,    0.99,    0.99,
  1.05,    1.05,    1.05,    1.05,
  0.33,    0.33,    0.33,    0.33,
  0.52,    0.52,    0.52,    0.52,
  0.37,    0.37,    0.37,    0.37,
  0.55,    0.55,    0.55,    0.55,
  1.27,    1.27,    1.27,    1.27,
  1.38,    1.38,    1.38,    1.38,
  1.19,    1.19,    1.19,    1.19,
  1.03,    1.03,    1.03,    1.03,
  0.19,    0.19,    0.19,    0.19,
  0.38,    0.38,    0.38,    0.38,
  0.72,    0.72,    0.72,    0.72,
  0.68,    0.68,    0.68,    0.68,
  1,       1,       1,       1,
  1.47,    1.47,    1.47,    1.47,
  1.8,     1.8,     1.8,     1.8,
  2.09,    2.09,    2.09,    2.09,
  2.46,    2.46,    2.46,    2.46,
  1.68,    1.68,    1.68,    1.68,
  2.63,    2.63,    2.63,    2.63,
  2.92,    2.92,    2.92,    2.92,
  2.7,     2.7,     2.7,     2.7,
  2.08,    2.08,    2.08,    2.08,
  2.34,    2.34,    2.34,    2.34,
  2.3,     2.3,     2.3,     2.3,
  2.35,    2.35,    2.35,    2.35,
  2.07,    2.07,    2.07,    2.07,
  2.22,    2.22,    2.22,    2.22,
  2.39,    2.39,    2.39,    2.39,
  2.43,    2.43,    2.43,    2.43,
  2.42,    2.42,    2.42,    2.42,
  2.64,    2.64,    2.64,    2.64,
  2.25,    2.25,    2.25,    2.25,
  2.58,    2.58,    2.58,    2.58,
  1.93,    1.93,    1.93,    1.93,
  0.99,    0.99,    0.99,    0.99,
  1.15,    1.15,    1.15,    1.15,
  2.17,    2.17,    2.17,    2.17,
  1.99,    1.99,    1.99,    1.99,
  1.22,    1.22,    1.22,    1.22,
  1.44,    1.44,    1.44,    1.44,
  1.38,    1.38,    1.38,    1.38,
  1.45,    1.45,    1.45,    1.45,
  1.53,    1.53,    1.53,    1.53,
  1.58,    1.58,    1.58,    1.58,
  1.74,    1.74,    1.74,    1.74,
  1.4,     1.4,     1.4,     1.4,
  2.23,    2.23,    2.23,    2.23,
  3.1,     3.1,     3.1,     3.1,
  3.19,    3.19,    3.19,    3.19,
  2.89,    2.89,    2.89,    2.89,
  3.07,    3.07,    3.07,    3.07,
  2.98,    2.98,    2.98,    2.98,
  3.16,    3.16,    3.16,    3.16,
  3.24,    3.24,    3.24,    3.24,
  3.38,    3.38,    3.38,    3.38,
  3.54,    3.54,    3.54,    3.54,
  3.81,    3.81,    3.81,    3.81,
  3.05,    3.05,    3.05,    3.05,
  3.64,    3.64,    3.64,    3.64,
  3.06,    3.06,    3.06,    3.06,
  3,       3,       3,       3,
  2.98,    2.98,    2.98,    2.98,
  2.59,    2.59,    2.59,    2.59,
  2.88,    2.88,    2.88,    2.88,
  2.68,    2.68,    2.68,    2.68,
  2.85,    2.85,    2.85,    2.85,
  2.9,     2.9,     2.9,     2.9,
  2.86,    2.86,    2.86,    2.86,
  3.58,    3.58,    3.58,    3.58,
  3.63,    3.63,    3.63,    3.63,
  3.22,    3.22,    3.22,    3.22,
  3.11,    3.11,    3.11,    3.11,
  2.64,    2.64,    2.64,    2.64,
  2.71,    2.71,    2.71,    2.71,
  2.67,    2.67,    2.67,    2.67,
  2.97,    2.97,    2.97,    2.97,
  2.7,     2.7,     2.7,     2.7,
  2.41,    2.41,    2.41,    2.41,
  2.01,    2.01,    2.01,    2.01,
  2.72,    2.72,    2.72,    2.72,
  2.68,    2.68,    2.68,    2.68,
  2.87,    2.87,    2.87,    2.87,
  3.21,    3.21,    3.21,    3.21,
  3.5,     3.5,     3.5,     3.5,
  2.86,    2.86,    2.86,    2.86,
  2.54,    2.54,    2.54,    2.54,
  3.17,    3.17,    3.17,    3.17,
  3.01,    3.01,    3.01,    3.01,
  3.82,    3.82,    3.82,    3.82,
  3.4,     3.4,     3.4,     3.4,
  3.82,    3.82,    3.82,    3.82,
  3.65,    3.65,    3.65,    3.65,
  4.38,    4.38,    4.38,    4.38,
  4.06,    4.06,    4.06,    4.06,
  4.13,    4.13,    4.13,    4.13,
  4.17,    4.17,    4.17,    4.17,
  4.55,    4.55,    4.55,    4.55,
  4.92,    4.92,    4.92,    4.92,
  4.59,    4.59,    4.59,    4.59,
  4.75,    4.75,    4.75,    4.75,
  4.83,    4.83,    4.83,    4.83,
  4.54,    4.54,    4.54,    4.54,
  5.08,    5.08,    5.08,    5.08,
  5.11,    5.11,    5.11,    5.11,
  4.87,    4.87,    4.87,    4.87,
  4.49,    4.49,    4.49,    4.49,
  4.8,     4.8,     4.8,     4.8,
  3.9,     3.9,     3.9,     3.9,
  3.7,     3.7,     3.7,     3.7,
  3.41,    3.41,    3.41,    3.41,
  2.87,    2.87,    2.87,    2.87,
  2.7,     2.7,     2.7,     2.7,
  2.78,    2.78,    2.78,    2.78,
  2.75,    2.75,    2.75,    2.75,
  2.89,    2.89,    2.89,    2.89,
  3.13,    3.13,    3.13,    3.13,
  3.56,    3.56,    3.56,    3.56,
  3.45,    3.45,    3.45,    3.45,
  3.09,    3.09,    3.09,    3.09,
  2.96,    2.96,    2.96,    2.96,
  3.01,    3.01,    3.01,    3.01,
  3.04,    3.04,    3.04,    3.04,
  2.77,    2.77,    2.77,    2.77,
  2.87,    2.87,    2.87,    2.87,
  2.49,    2.49,    2.49,    2.49,
  2.35,    2.35,    2.35,    2.35,
  2.47,    2.47,    2.47,    2.47,
  2.61,    2.61,    2.61,    2.61,
  2.24,    2.24,    2.24,    2.24,
  2.44,    2.44,    2.44,    2.44,
  2.77,    2.77,    2.77,    2.77,
  1.98,    1.98,    1.98,    1.98,
  1.61,    1.61,    1.61,    1.61,
  2.11,    2.11,    2.11,    2.11,
  2.08,    2.08,    2.08,    2.08,
  2.24,    2.24,    2.24,    2.24,
  3.05,    3.05,    3.05,    3.05,
  2.56,    2.56,    2.56,    2.56,
  2.31,    2.31,    2.31,    2.31,
  2.24,    2.24,    2.24,    2.24,
  2.15,    2.15,    2.15,    2.15,
  2.54,    2.54,    2.54,    2.54,
  2.55,    2.55,    2.55,    2.55,
  3.2,     3.2,     3.2,     3.2,
  3.17,    3.17,    3.17,    3.17,
  2.67,    2.67,    2.67,    2.67,
  2.35,    2.35,    2.35,    2.35,
  2.68,    2.68,    2.68,    2.68,
  2.1,     2.1,     2.1,     2.1,
  2.11,    2.11,    2.11,    2.11,
  2.55,    2.55,    2.55,    2.55,
  2.49,    2.49,    2.49,    2.49,
  2.05,    2.05,    2.05,    2.05,
  2.18,    2.18,    2.18,    2.18,
  2.2,     2.2,     2.2,     2.2,
  2.4,     2.4,     2.4,     2.4,
  2.62,    2.62,    2.62,    2.62,
  2.03,    2.03,    2.03,    2.03,
  1.83,    1.83,    1.83,    1.83,
  2.43,    2.43,    2.43,    2.43,
  2.71,    2.71,    2.71,    2.71,
  2.86,    2.86,    2.86,    2.86,
  2.82,    2.82,    2.82,    2.82,
  2.81,    2.81,    2.81,    2.81,
  2.98,    2.98,    2.98,    2.98,
  3.13,    3.13,    3.13,    3.13,
  3.33,    3.33,    3.33,    3.33,
  2.77,    2.77,    2.77,    2.77,
  2.6,     2.6,     2.6,     2.6,
  2.24,    2.24,    2.24,    2.24,
  2.37,    2.37,    2.37,    2.37,
  2.41,    2.41,    2.41,    2.41,
  2.33,    2.33,    2.33,    2.33,
  2.49,    2.49,    2.49,    2.49,
  1.9,     1.9,     1.9,     1.9,
  1.18,    1.18,    1.18,    1.18,
  1.3,     1.3,     1.3,     1.3,
  2.27,    2.27,    2.27,    2.27,
  2.27,    2.27,    2.27,    2.27,
  2.37,    2.37,    2.37,    2.37,
  1.96,    1.96,    1.96,    1.96,
  1.32,    1.32,    1.32,    1.32,
  1.29,    1.29,    1.29,    1.29,
  1.26,    1.26,    1.26,    1.26,
  0.91,    0.91,    0.91,    0.91,
  0.92,    0.92,    0.92,    0.92,
  0.78,    0.78,    0.78,    0.78,
  0.58,    0.58,    0.58,    0.58,
  1.31,    1.31,    1.31,    1.31,
  1.85,    1.85,    1.85,    1.85,
  2.7,     2.7,     2.7,     2.7,
  2.94,    2.94,    2.94,    2.94,
  2.7,     2.7,     2.7,     2.7,
  3.15,    3.15,    3.15,    3.15,
  3.18,    3.18,    3.18,    3.18,
  2.33,    2.33,    2.33,    2.33,
  2,       2,       2,       2,
  3.25,    3.25,    3.25,    3.25,
  2.25,    2.25,    2.25,    2.25,
  2.5,     2.5,     2.5,     2.5,
  2.6,     2.6,     2.6,     2.6,
  2.33,    2.33,    2.33,    2.33,
  2.63,    2.63,    2.63,    2.63,
  2.03,    2.03,    2.03,    2.03,
  1.33,    1.33,    1.33,    1.33,
  1.91,    1.91,    1.91,    1.91,
  3.09,    3.09,    3.09,    3.09,
  2.65,    2.65,    2.65,    2.65,
  2.3,     2.3,     2.3,     2.3,
  2.41,    2.41,    2.41,    2.41,
  2.29,    2.29,    2.29,    2.29,
  2.46,    2.46,    2.46,    2.46,
  2.74,    2.74,    2.74,    2.74,
  2.47,    2.47,    2.47,    2.47,
  1.34,    1.34,    1.34,    1.34,
  1.8,     1.8,     1.8,     1.8,
  1.89,    1.89,    1.89,    1.89,
  1.7,     1.7,     1.7,     1.7,
  2.07,    2.07,    2.07,    2.07,
  2.01,    2.01,    2.01,    2.01,
  1.95,    1.95,    1.95,    1.95,
  2.02,    2.02,    2.02,    2.02,
  1.97,    1.97,    1.97,    1.97,
  2.12,    2.12,    2.12,    2.12,
  1.91,    1.91,    1.91,    1.91,
  1.85,    1.85,    1.85,    1.85,
  1.74,    1.74,    1.74,    1.74,
  1.91,    1.91,    1.91,    1.91,
  2.3,     2.3,     2.3,     2.3,
  2.28,    2.28,    2.28,    2.28,
  2.4,     2.4,     2.4,     2.4,
  1.84,    1.84,    1.84,    1.84,
  2.63,    2.63,    2.63,    2.63,
  2.01,    2.01,    2.01,    2.01,
  2.01,    2.01,    2.01,    2.01,
  2.65,    2.65,    2.65,    2.65,
  2.87,    2.87,    2.87,    2.87,
  4.19,    4.19,    4.19,    4.19,
  3.12,    3.12,    3.12,    3.12,
  3.46,    3.46,    3.46,    3.46,
  3.39,    3.39,    3.39,    3.39,
  3.37,    3.37,    3.37,    3.37,
  3.35,    3.35,    3.35,    3.35,
  3.73,    3.73,    3.73,    3.73,
  3.62,    3.62,    3.62,    3.62,
  3.8,     3.8,     3.8,     3.8,
  3.42,    3.42,    3.42,    3.42,
  3.78,    3.78,    3.78,    3.78,
  3.74,    3.74,    3.74,    3.74,
  3.37,    3.37,    3.37,    3.37,
  2.91,    2.91,    2.91,    2.91,
  3.17,    3.17,    3.17,    3.17,
  2.18,    2.18,    2.18,    2.18,
  2.31,    2.31,    2.31,    2.31,
  2.51,    2.51,    2.51,    2.51,
  2.57,    2.57,    2.57,    2.57,
  2,       2,       2,       2,
  1.95,    1.95,    1.95,    1.95,
  2.43,    2.43,    2.43,    2.43,
  1.94,    1.94,    1.94,    1.94,
  2.26,    2.26,    2.26,    2.26,
  2.09,    2.09,    2.09,    2.09,
  1.92,    1.92,    1.92,    1.92,
  2.01,    2.01,    2.01,    2.01,
  1.31,    1.31,    1.31,    1.31,
  1.14,    1.14,    1.14,    1.14,
  1.12,    1.12,    1.12,    1.12,
  1.84,    1.84,    1.84,    1.84,
  1.67,    1.67,    1.67,    1.67,
  1.85,    1.85,    1.85,    1.85,
  1.53,    1.53,    1.53,    1.53,
  1.48,    1.48,    1.48,    1.48,
  1.59,    1.59,    1.59,    1.59,
  1.51,    1.51,    1.51,    1.51,
  1.72,    1.72,    1.72,    1.72,
  1.38,    1.38,    1.38,    1.38,
  0.96,    0.96,    0.96,    0.96,
  1.16,    1.16,    1.16,    1.16,
  1.58,    1.58,    1.58,    1.58,
  1.93,    1.93,    1.93,    1.93,
  1.98,    1.98,    1.98,    1.98,
  2.12,    2.12,    2.12,    2.12,
  1.83,    1.83,    1.83,    1.83,
  2.7,     2.7,     2.7,     2.7,
  3.23,    3.23,    3.23,    3.23,
  2.85,    2.85,    2.85,    2.85,
  2.55,    2.55,    2.55,    2.55,
  3.17,    3.17,    3.17,    3.17,
  2.96,    2.96,    2.96,    2.96,
  2.98,    2.98,    2.98,    2.98,
  2.91,    2.91,    2.91,    2.91,
  3.22,    3.22,    3.22,    3.22,
  2.9,     2.9,     2.9,     2.9,
  3.22,    3.22,    3.22,    3.22,
  3.28,    3.28,    3.28,    3.28,
  2.88,    2.88,    2.88,    2.88,
  3.04,    3.04,    3.04,    3.04,
  3.75,    3.75,    3.75,    3.75,
  2.78,    2.78,    2.78,    2.78,
  3.09,    3.09,    3.09,    3.09,
  2.59,    2.59,    2.59,    2.59,
  1.98,    1.98,    1.98,    1.98,
  1.81,    1.81,    1.81,    1.81,
  1.51,    1.51,    1.51,    1.51,
  1.86,    1.86,    1.86,    1.86,
  2.28,    2.28,    2.28,    2.28,
  1.97,    1.97,    1.97,    1.97,
  1.42,    1.42,    1.42,    1.42,
  1.58,    1.58,    1.58,    1.58,
  1.86,    1.86,    1.86,    1.86,
  2.09,    2.09,    2.09,    2.09,
  1.59,    1.59,    1.59,    1.59,
  1.53,    1.53,    1.53,    1.53,
  1.4,     1.4,     1.4,     1.4,
  0.42,    0.42,    0.42,    0.42,
  1.21,    1.21,    1.21,    1.21,
  1.64,    1.64,    1.64,    1.64,
  1.97,    1.97,    1.97,    1.97,
  1.63,    1.63,    1.63,    1.63,
  1.85,    1.85,    1.85,    1.85,
  2.27,    2.27,    2.27,    2.27,
  1.78,    1.78,    1.78,    1.78,
  1.65,    1.65,    1.65,    1.65,
  1.48,    1.48,    1.48,    1.48,
  2.16,    2.16,    2.16,    2.16,
  1.24,    1.24,    1.24,    1.24,
  0.78,    0.78,    0.78,    0.78,
  0.96,    0.96,    0.96,    0.96,
  1.43,    1.43,    1.43,    1.43,
  2.2,     2.2,     2.2,     2.2,
  1.59,    1.59,    1.59,    1.59,
  1.34,    1.34,    1.34,    1.34,
  1.46,    1.46,    1.46,    1.46,
  1.9,     1.9,     1.9,     1.9,
  2.07,    2.07,    2.07,    2.07,
  1.92,    1.92,    1.92,    1.92,
  1.87,    1.87,    1.87,    1.87,
  1.9,     1.9,     1.9,     1.9,
  1.99,    1.99,    1.99,    1.99,
  1.11,    1.11,    1.11,    1.11,
  0.79,    0.79,    0.79,    0.79,
  1.64,    1.64,    1.64,    1.64,
  1.59,    1.59,    1.59,    1.59,
  2.19,    2.19,    2.19,    2.19,
  1.43,    1.43,    1.43,    1.43,
  1.57,    1.57,    1.57,    1.57,
  2.19,    2.19,    2.19,    2.19,
  1.92,    1.92,    1.92,    1.92,
  1.98,    1.98,    1.98,    1.98,
  1.87,    1.87,    1.87,    1.87,
  1.94,    1.94,    1.94,    1.94,
  2.28,    2.28,    2.28,    2.28,
  2.13,    2.13,    2.13,    2.13,
  2.27,    2.27,    2.27,    2.27,
  2.28,    2.28,    2.28,    2.28,
  2.09,    2.09,    2.09,    2.09,
  2.24,    2.24,    2.24,    2.24,
  2.52,    2.52,    2.52,    2.52,
  2.25,    2.25,    2.25,    2.25,
  2.34,    2.34,    2.34,    2.34,
  2.39,    2.39,    2.39,    2.39,
  2,       2,       2,       2,
  1.95,    1.95,    1.95,    1.95,
  1.96,    1.96,    1.96,    1.96,
  1.94,    1.94,    1.94,    1.94,
  1.73,    1.73,    1.73,    1.73,
  1.68,    1.68,    1.68,    1.68,
  1.55,    1.55,    1.55,    1.55,
  1.81,    1.81,    1.81,    1.81,
  1.46,    1.46,    1.46,    1.46,
  1.58,    1.58,    1.58,    1.58,
  1.59,    1.59,    1.59,    1.59,
  1.52,    1.52,    1.52,    1.52,
  1.4,     1.4,     1.4,     1.4,
  1.6,     1.6,     1.6,     1.6,
  1.47,    1.47,    1.47,    1.47,
  0.81,    0.81,    0.81,    0.81,
  0.45,    0.45,    0.45,    0.45,
  0.58,    0.58,    0.58,    0.58,
  0.5,     0.5,     0.5,     0.5,
  0.43,    0.43,    0.43,    0.43,
  0.98,    0.98,    0.98,    0.98,
  1.07,    1.07,    1.07,    1.07,
  1.22,    1.22,    1.22,    1.22,
  1.93,    1.93,    1.93,    1.93,
  1.42,    1.42,    1.42,    1.42,
  1.91,    1.91,    1.91,    1.91,
  1.81,    1.81,    1.81,    1.81,
  1.91,    1.91,    1.91,    1.91,
  1.55,    1.55,    1.55,    1.55,
  1.47,    1.47,    1.47,    1.47,
  1.29,    1.29,    1.29,    1.29,
  2.24,    2.24,    2.24,    2.24,
  1.42,    1.42,    1.42,    1.42,
  2.95,    2.95,    2.95,    2.95,
  2.52,    2.52,    2.52,    2.52,
  1.96,    1.96,    1.96,    1.96,
  1.9,     1.9,     1.9,     1.9,
  1.63,    1.63,    1.63,    1.63,
  1.78,    1.78,    1.78,    1.78,
  1.9,     1.9,     1.9,     1.9,
  1.78,    1.78,    1.78,    1.78,
  2.18,    2.18,    2.18,    2.18,
  1.61,    1.61,    1.61,    1.61,
  1.63,    1.63,    1.63,    1.63,
  1.87,    1.87,    1.87,    1.87,
  1.32,    1.32,    1.32,    1.32,
  2,       2,       2,       2,
  2.61,    2.61,    2.61,    2.61,
  0.84,    0.84,    0.84,    0.84,
  0.74,    0.74,    0.74,    0.74,
  1.71,    1.71,    1.71,    1.71,
  2.72,    2.72,    2.72,    2.72,
  1.49,    1.49,    1.49,    1.49,
  0.12,    0.12,    0.12,    0.12,
  1.16,    1.16,    1.16,    1.16,
  2.48,    2.48,    2.48,    2.48,
  2.62,    2.62,    2.62,    2.62,
  1.34,    1.34,    1.34,    1.34,
  1.75,    1.75,    1.75,    1.75,
  2.11,    2.11,    2.11,    2.11,
  1.47,    1.47,    1.47,    1.47,
  1.62,    1.62,    1.62,    1.62,
  0.95,    0.95,    0.95,    0.95,
  1.32,    1.32,    1.32,    1.32,
  0.88,    0.88,    0.88,    0.88,
  1.67,    1.67,    1.67,    1.67,
  2.78,    2.78,    2.78,    2.78,
  2.47,    2.47,    2.47,    2.47,
  2.91,    2.91,    2.91,    2.91,
  2.78,    2.78,    2.78,    2.78,
  3.03,    3.03,    3.03,    3.03,
  2.77,    2.77,    2.77,    2.77,
  2.57,    2.57,    2.57,    2.57,
  2.56,    2.56,    2.56,    2.56,
  2.41,    2.41,    2.41,    2.41,
  3.34,    3.34,    3.34,    3.34,
  2.67,    2.67,    2.67,    2.67,
  2.73,    2.73,    2.73,    2.73,
  2.3,     2.3,     2.3,     2.3,
  2.69,    2.69,    2.69,    2.69,
  3.08,    3.08,    3.08,    3.08,
  2.31,    2.31,    2.31,    2.31,
  1.75,    1.75,    1.75,    1.75,
  2.1,     2.1,     2.1,     2.1,
  1.4,     1.4,     1.4,     1.4,
  1.61,    1.61,    1.61,    1.61,
  1.66,    1.66,    1.66,    1.66,
  1.93,    1.93,    1.93,    1.93,
  1.93,    1.93,    1.93,    1.93,
  2.48,    2.48,    2.48,    2.48,
  2.49,    2.49,    2.49,    2.49,
  3.07,    3.07,    3.07,    3.07,
  3,       3,       3,       3,
  2.73,    2.73,    2.73,    2.73,
  2.78,    2.78,    2.78,    2.78,
  2.79,    2.79,    2.79,    2.79,
  2.86,    2.86,    2.86,    2.86,
  2.94,    2.94,    2.94,    2.94,
  2.83,    2.83,    2.83,    2.83,
  2.56,    2.56,    2.56,    2.56,
  2.46,    2.46,    2.46,    2.46,
  2.74,    2.74,    2.74,    2.74,
  3.19,    3.19,    3.19,    3.19,
  3,       3,       3,       3,
  2.66,    2.66,    2.66,    2.66,
  3.38,    3.38,    3.38,    3.38,
  3.01,    3.01,    3.01,    3.01,
  2.59,    2.59,    2.59,    2.59,
  1.89,    1.89,    1.89,    1.89,
  1.04,    1.04,    1.04,    1.04,
  1.98,    1.98,    1.98,    1.98,
  2.65,    2.65,    2.65,    2.65,
  2.56,    2.56,    2.56,    2.56,
  3.51,    3.51,    3.51,    3.51,
  3.97,    3.97,    3.97,    3.97,
  3.02,    3.02,    3.02,    3.02,
  3.58,    3.58,    3.58,    3.58,
  3.59,    3.59,    3.59,    3.59,
  4.07,    4.07,    4.07,    4.07,
  3.98,    3.98,    3.98,    3.98,
  3.74,    3.74,    3.74,    3.74,
  4.18,    4.18,    4.18,    4.18,
  3.8,     3.8,     3.8,     3.8,
  3.17,    3.17,    3.17,    3.17,
  3.25,    3.25,    3.25,    3.25,
  3.64,    3.64,    3.64,    3.64,
  3.63,    3.63,    3.63,    3.63,
  4.06,    4.06,    4.06,    4.06,
  4.02,    4.02,    4.02,    4.02,
  3.76,    3.76,    3.76,    3.76,
  4.58,    4.58,    4.58,    4.58,
  4.21,    4.21,    4.21,    4.21,
  3.71,    3.71,    3.71,    3.71,
  3.62,    3.62,    3.62,    3.62,
  2.38,    2.38,    2.38,    2.38,
  2.77,    2.77,    2.77,    2.77,
  2.82,    2.82,    2.82,    2.82,
  2.07,    2.07,    2.07,    2.07,
  1.85,    1.85,    1.85,    1.85,
  1.67,    1.67,    1.67,    1.67,
  1.75,    1.75,    1.75,    1.75,
  1.45,    1.45,    1.45,    1.45,
  1.76,    1.76,    1.76,    1.76,
  1.55,    1.55,    1.55,    1.55,
  1.58,    1.58,    1.58,    1.58,
  1.5,     1.5,     1.5,     1.5,
  2.12,    2.12,    2.12,    2.12,
  1.92,    1.92,    1.92,    1.92,
  1.9,     1.9,     1.9,     1.9,
  0.95,    0.95,    0.95,    0.95,
  1.03,    1.03,    1.03,    1.03,
  0.72,    0.72,    0.72,    0.72,
  1.02,    1.02,    1.02,    1.02,
  1.75,    1.75,    1.75,    1.75,
  1.06,    1.06,    1.06,    1.06,
  1.33,    1.33,    1.33,    1.33,
  1.94,    1.94,    1.94,    1.94,
  1.63,    1.63,    1.63,    1.63,
  1.96,    1.96,    1.96,    1.96,
  1.82,    1.82,    1.82,    1.82,
  1.77,    1.77,    1.77,    1.77,
  2.24,    2.24,    2.24,    2.24,
  3.27,    3.27,    3.27,    3.27,
  3.52,    3.52,    3.52,    3.52,
  4.13,    4.13,    4.13,    4.13,
  3.87,    3.87,    3.87,    3.87,
  4.23,    4.23,    4.23,    4.23,
  3.56,    3.56,    3.56,    3.56,
  3.01,    3.01,    3.01,    3.01,
  3.1,     3.1,     3.1,     3.1,
  3.02,    3.02,    3.02,    3.02,
  3.2,     3.2,     3.2,     3.2,
  2.49,    2.49,    2.49,    2.49,
  2.09,    2.09,    2.09,    2.09,
  2.53,    2.53,    2.53,    2.53,
  2.06,    2.06,    2.06,    2.06,
  2.62,    2.62,    2.62,    2.62,
  2.69,    2.69,    2.69,    2.69,
  1.76,    1.76,    1.76,    1.76,
  1.45,    1.45,    1.45,    1.45,
  1.3,     1.3,     1.3,     1.3,
  0.69,    0.69,    0.69,    0.69,
  1.83,    1.83,    1.83,    1.83,
  1.81,    1.81,    1.81,    1.81,
  2,       2,       2,       2,
  2.04,    2.04,    2.04,    2.04,
  2,       2,       2,       2,
  1.68,    1.68,    1.68,    1.68,
  0.96,    0.96,    0.96,    0.96,
  0.91,    0.91,    0.91,    0.91,
  1.11,    1.11,    1.11,    1.11,
  1.64,    1.64,    1.64,    1.64,
  1.55,    1.55,    1.55,    1.55,
  1.75,    1.75,    1.75,    1.75,
  1.8,     1.8,     1.8,     1.8,
  1.63,    1.63,    1.63,    1.63,
  1.96,    1.96,    1.96,    1.96,
  2.03,    2.03,    2.03,    2.03,
  2.24,    2.24,    2.24,    2.24,
  2.2,     2.2,     2.2,     2.2,
  2.17,    2.17,    2.17,    2.17,
  2.22,    2.22,    2.22,    2.22,
  2.12,    2.12,    2.12,    2.12,
  1.94,    1.94,    1.94,    1.94,
  1.71,    1.71,    1.71,    1.71,
  1.71,    1.71,    1.71,    1.71,
  1.36,    1.36,    1.36,    1.36,
  1.23,    1.23,    1.23,    1.23,
  1.75,    1.75,    1.75,    1.75,
  2.21,    2.21,    2.21,    2.21,
  1.77,    1.77,    1.77,    1.77,
  2.15,    2.15,    2.15,    2.15,
  2.29,    2.29,    2.29,    2.29,
  2.06,    2.06,    2.06,    2.06,
  2.3,     2.3,     2.3,     2.3,
  2.3,     2.3,     2.3,     2.3,
  2.88,    2.88,    2.88,    2.88,
  2.61,    2.61,    2.61,    2.61,
  2.22,    2.22,    2.22,    2.22,
  2.04,    2.04,    2.04,    2.04,
  2.03,    2.03,    2.03,    2.03,
  2.29,    2.29,    2.29,    2.29,
  1.83,    1.83,    1.83,    1.83,
  2.19,    2.19,    2.19,    2.19,
  2.23,    2.23,    2.23,    2.23,
  1.97,    1.97,    1.97,    1.97,
  1.56,    1.56,    1.56,    1.56,
  1.55,    1.55,    1.55,    1.55,
  1.3,     1.3,     1.3,     1.3,
  1.91,    1.91,    1.91,    1.91,
  1.59,    1.59,    1.59,    1.59,
  1.82,    1.82,    1.82,    1.82,
  2.06,    2.06,    2.06,    2.06,
  2.14,    2.14,    2.14,    2.14,
  2.24,    2.24,    2.24,    2.24,
  2.09,    2.09,    2.09,    2.09,
  2.21,    2.21,    2.21,    2.21,
  2.21,    2.21,    2.21,    2.21,
  2.33,    2.33,    2.33,    2.33,
  2.45,    2.45,    2.45,    2.45,
  2.37,    2.37,    2.37,    2.37,
  2.24,    2.24,    2.24,    2.24,
  1.6,     1.6,     1.6,     1.6,
  1.73,    1.73,    1.73,    1.73,
  1.9,     1.9,     1.9,     1.9,
  1.88,    1.88,    1.88,    1.88,
  1.84,    1.84,    1.84,    1.84,
  1.75,    1.75,    1.75,    1.75,
  1.74,    1.74,    1.74,    1.74,
  1.57,    1.57,    1.57,    1.57,
  1.42,    1.42,    1.42,    1.42,
  1.47,    1.47,    1.47,    1.47,
  1.73,    1.73,    1.73,    1.73,
  1.69,    1.69,    1.69,    1.69,
  2.24,    2.24,    2.24,    2.24,
  1.88,    1.88,    1.88,    1.88,
  2.35,    2.35,    2.35,    2.35,
  1.98,    1.98,    1.98,    1.98,
  1.7,     1.7,     1.7,     1.7,
  2.03,    2.03,    2.03,    2.03,
  2.6,     2.6,     2.6,     2.6,
  2.28,    2.28,    2.28,    2.28,
  2.37,    2.37,    2.37,    2.37,
  2.65,    2.65,    2.65,    2.65,
  2.23,    2.23,    2.23,    2.23,
  2.39,    2.39,    2.39,    2.39,
  2.7,     2.7,     2.7,     2.7,
  2.7,     2.7,     2.7,     2.7,
  2.24,    2.24,    2.24,    2.24,
  1.82,    1.82,    1.82,    1.82,
  2.31,    2.31,    2.31,    2.31,
  2.13,    2.13,    2.13,    2.13,
  1.99,    1.99,    1.99,    1.99,
  1.81,    1.81,    1.81,    1.81,
  1.65,    1.65,    1.65,    1.65,
  1.83,    1.83,    1.83,    1.83,
  1.7,     1.7,     1.7,     1.7,
  1.43,    1.43,    1.43,    1.43,
  1.13,    1.13,    1.13,    1.13,
  1.11,    1.11,    1.11,    1.11,
  1.37,    1.37,    1.37,    1.37,
  1.09,    1.09,    1.09,    1.09,
  1.15,    1.15,    1.15,    1.15,
  1.09,    1.09,    1.09,    1.09,
  1.04,    1.04,    1.04,    1.04,
  1.02,    1.02,    1.02,    1.02,
  1.06,    1.06,    1.06,    1.06,
  1.06,    1.06,    1.06,    1.06,
  0.94,    0.94,    0.94,    0.94,
  0.73,    0.73,    0.73,    0.73,
  1.04,    1.04,    1.04,    1.04,
  0.32,    0.32,    0.32,    0.32,
  0.26,    0.26,    0.26,    0.26,
  0.74,    0.74,    0.74,    0.74,
  0.9,     0.9,     0.9,     0.9,
  0.77,    0.77,    0.77,    0.77,
  1.31,    1.31,    1.31,    1.31,
  0.23,    0.23,    0.23,    0.23,
  0.28,    0.28,    0.28,    0.28,
  0.47,    0.47,    0.47,    0.47,
  0.22,    0.22,    0.22,    0.22,
  0.22,    0.22,    0.22,    0.22,
  0.56,    0.56,    0.56,    0.56,
  0.36,    0.36,    0.36,    0.36,
  1.07,    1.07,    1.07,    1.07,
  1.03,    1.03,    1.03,    1.03,
  0.36,    0.36,    0.36,    0.36,
  0.76,    0.76,    0.76,    0.76,
  0.78,    0.78,    0.78,    0.78,
  0.76,    0.76,    0.76,    0.76,
  1.51,    1.51,    1.51,    1.51,
  1.91,    1.91,    1.91,    1.91,
  2.43,    2.43,    2.43,    2.43,
  2.14,    2.14,    2.14,    2.14,
  2.02,    2.02,    2.02,    2.02,
  2.07,    2.07,    2.07,    2.07,
  1.93,    1.93,    1.93,    1.93,
  2.52,    2.52,    2.52,    2.52,
  2.12,    2.12,    2.12,    2.12,
  2.28,    2.28,    2.28,    2.28,
  1.79,    1.79,    1.79,    1.79,
  1.47,    1.47,    1.47,    1.47,
  1.14,    1.14,    1.14,    1.14,
  1.25,    1.25,    1.25,    1.25,
  1.29,    1.29,    1.29,    1.29,
  1.66,    1.66,    1.66,    1.66,
  1.74,    1.74,    1.74,    1.74,
  2.2,     2.2,     2.2,     2.2,
  2.07,    2.07,    2.07,    2.07,
  2.08,    2.08,    2.08,    2.08,
  2.04,    2.04,    2.04,    2.04,
  2.07,    2.07,    2.07,    2.07,
  2.3,     2.3,     2.3,     2.3,
  2.55,    2.55,    2.55,    2.55,
  2.58,    2.58,    2.58,    2.58,
  2.59,    2.59,    2.59,    2.59,
  2.63,    2.63,    2.63,    2.63,
  2.41,    2.41,    2.41,    2.41,
  2.63,    2.63,    2.63,    2.63,
  2.58,    2.58,    2.58,    2.58,
  2.45,    2.45,    2.45,    2.45,
  2.3,     2.3,     2.3,     2.3,
  2.38,    2.38,    2.38,    2.38,
  2.54,    2.54,    2.54,    2.54,
  2.38,    2.38,    2.38,    2.38,
  2.41,    2.41,    2.41,    2.41,
  2.15,    2.15,    2.15,    2.15,
  1.82,    1.82,    1.82,    1.82,
  1.76,    1.76,    1.76,    1.76,
  2.01,    2.01,    2.01,    2.01,
  2.05,    2.05,    2.05,    2.05,
  2.43,    2.43,    2.43,    2.43,
  1.67,    1.67,    1.67,    1.67,
  1.58,    1.58,    1.58,    1.58,
  1.68,    1.68,    1.68,    1.68,
  1.84,    1.84,    1.84,    1.84,
  2.33,    2.33,    2.33,    2.33,
  2.5,     2.5,     2.5,     2.5,
  2.39,    2.39,    2.39,    2.39,
  2.42,    2.42,    2.42,    2.42,
  2.91,    2.91,    2.91,    2.91,
  2.59,    2.59,    2.59,    2.59,
  2.46,    2.46,    2.46,    2.46,
  2.73,    2.73,    2.73,    2.73,
  2.74,    2.74,    2.74,    2.74,
  2.49,    2.49,    2.49,    2.49,
  2.29,    2.29,    2.29,    2.29,
  1.99,    1.99,    1.99,    1.99,
  1.96,    1.96,    1.96,    1.96,
  2.06,    2.06,    2.06,    2.06,
  1.74,    1.74,    1.74,    1.74,
  0.64,    0.64,    0.64,    0.64,
  0.81,    0.81,    0.81,    0.81,
  1.18,    1.18,    1.18,    1.18,
  1.69,    1.69,    1.69,    1.69,
  2.16,    2.16,    2.16,    2.16,
  2.07,    2.07,    2.07,    2.07,
  2.71,    2.71,    2.71,    2.71,
  2.74,    2.74,    2.74,    2.74,
  2.72,    2.72,    2.72,    2.72,
  2.76,    2.76,    2.76,    2.76,
  3.21,    3.21,    3.21,    3.21,
  2.79,    2.79,    2.79,    2.79,
  2.052,   2.052,   2.052,   2.052,
  1.777,   1.777,   1.777,   1.777,
  1.666,   1.666,   1.666,   1.666,
  1.924,   1.924,   1.924,   1.924,
  1.887,   1.887,   1.887,   1.887,
  1.824,   1.824,   1.824,   1.824,
  1.587,   1.587,   1.587,   1.587,
  1.711,   1.711,   1.711,   1.711,
  2,       2,       2,       2,
  1.9,     1.9,     1.9,     1.9,
  1.64,    1.64,    1.64,    1.64,
  1.38,    1.38,    1.38,    1.38,
  1.05,    1.05,    1.05,    1.05,
  0.57,    0.57,    0.57,    0.57,
  0.54,    0.54,    0.54,    0.54,
  1.23,    1.23,    1.23,    1.23,
  1.21,    1.21,    1.21,    1.21,
  1.5,     1.5,     1.5,     1.5,
  1.65,    1.65,    1.65,    1.65,
  1.35,    1.35,    1.35,    1.35,
  1.22,    1.22,    1.22,    1.22,
  0.9,     0.9,     0.9,     0.9,
  0.29,    0.29,    0.29,    0.29,
  0.96,    0.96,    0.96,    0.96,
  1.19,    1.19,    1.19,    1.19,
  2.37,    2.37,    2.37,    2.37,
  2.76,    2.76,    2.76,    2.76,
  3.86,    3.86,    3.86,    3.86,
  3.97,    3.97,    3.97,    3.97,
  3.45,    3.45,    3.45,    3.45,
  2.18,    2.18,    2.18,    2.18,
  1.16,    1.16,    1.16,    1.16,
  6.21,    6.21,    6.21,    6.21,
  2.28,    2.28,    2.28,    2.28,
  1.87,    1.87,    1.87,    1.87,
  1.97,    1.97,    1.97,    1.97,
  0.61,    0.61,    0.61,    0.61,
  1.04,    1.04,    1.04,    1.04,
  1.19,    1.19,    1.19,    1.19,
  0.91,    0.91,    0.91,    0.91,
  0.39,    0.39,    0.39,    0.39,
  0.71,    0.71,    0.71,    0.71,
  1.16,    1.16,    1.16,    1.16,
  1.69,    1.69,    1.69,    1.69,
  1.94,    1.94,    1.94,    1.94,
  1.62,    1.62,    1.62,    1.62,
  2.44,    2.44,    2.44,    2.44,
  2.18,    2.18,    2.18,    2.18,
  2.27,    2.27,    2.27,    2.27,
  1.85,    1.85,    1.85,    1.85,
  1.42,    1.42,    1.42,    1.42,
  1.85,    1.85,    1.85,    1.85,
  1.54,    1.54,    1.54,    1.54,
  1.23,    1.23,    1.23,    1.23,
  1.16,    1.16,    1.16,    1.16,
  1.32,    1.32,    1.32,    1.32,
  1.23,    1.23,    1.23,    1.23,
  1.29,    1.29,    1.29,    1.29,
  1.51,    1.51,    1.51,    1.51,
  1.12,    1.12,    1.12,    1.12,
  1.23,    1.23,    1.23,    1.23,
  1.56,    1.56,    1.56,    1.56,
  1.14,    1.14,    1.14,    1.14,
  0.8,     0.8,     0.8,     0.8,
  1.05,    1.05,    1.05,    1.05,
  1.04,    1.04,    1.04,    1.04,
  0.8,     0.8,     0.8,     0.8,
  1.14,    1.14,    1.14,    1.14,
  0.96,    0.96,    0.96,    0.96,
  0.8,     0.8,     0.8,     0.8,
  1.08,    1.08,    1.08,    1.08,
  1.01,    1.01,    1.01,    1.01,
  0.9,     0.9,     0.9,     0.9,
  0.53,    0.53,    0.53,    0.53,
  0.83,    0.83,    0.83,    0.83,
  0.96,    0.96,    0.96,    0.96,
  1.49,    1.49,    1.49,    1.49,
  1.53,    1.53,    1.53,    1.53,
  1.59,    1.59,    1.59,    1.59,
  1.63,    1.63,    1.63,    1.63,
  2.15,    2.15,    2.15,    2.15,
  1.09,    1.09,    1.09,    1.09,
  1.34,    1.34,    1.34,    1.34,
  1.35,    1.35,    1.35,    1.35,
  1.73,    1.73,    1.73,    1.73,
  1.72,    1.72,    1.72,    1.72,
  1.47,    1.47,    1.47,    1.47,
  1.62,    1.62,    1.62,    1.62,
  1.12,    1.12,    1.12,    1.12,
  0.48,    0.48,    0.48,    0.48,
  0.45,    0.45,    0.45,    0.45,
  0.98,    0.98,    0.98,    0.98,
  0.85,    0.85,    0.85,    0.85,
  1.15,    1.15,    1.15,    1.15,
  1.13,    1.13,    1.13,    1.13,
  1.91,    1.91,    1.91,    1.91,
  2.33,    2.33,    2.33,    2.33,
  1.98,    1.98,    1.98,    1.98,
  2.35,    2.35,    2.35,    2.35,
  2.4,     2.4,     2.4,     2.4,
  1.78,    1.78,    1.78,    1.78,
  1.89,    1.89,    1.89,    1.89,
  1.64,    1.64,    1.64,    1.64,
  1.75,    1.75,    1.75,    1.75,
  1.02,    1.02,    1.02,    1.02,
  1.08,    1.08,    1.08,    1.08,
  1.42,    1.42,    1.42,    1.42,
  1.67,    1.67,    1.67,    1.67,
  1.52,    1.52,    1.52,    1.52,
  1.25,    1.25,    1.25,    1.25,
  1.62,    1.62,    1.62,    1.62,
  1.88,    1.88,    1.88,    1.88,
  1.78,    1.78,    1.78,    1.78,
  2.09,    2.09,    2.09,    2.09,
  1.84,    1.84,    1.84,    1.84,
  2.57,    2.57,    2.57,    2.57,
  2.11,    2.11,    2.11,    2.11,
  2.19,    2.19,    2.19,    2.19,
  3.11,    3.11,    3.11,    3.11,
  2.81,    2.81,    2.81,    2.81,
  3.08,    3.08,    3.08,    3.08,
  3.06,    3.06,    3.06,    3.06,
  2.84,    2.84,    2.84,    2.84,
  3.2,     3.2,     3.2,     3.2,
  2.81,    2.81,    2.81,    2.81,
  3.58,    3.58,    3.58,    3.58,
  2.54,    2.54,    2.54,    2.54,
  2.56,    2.56,    2.56,    2.56,
  2.96,    2.96,    2.96,    2.96,
  0.84,    0.84,    0.84,    0.84,
  0.98,    0.98,    0.98,    0.98,
  1.25,    1.25,    1.25,    1.25,
  1.85,    1.85,    1.85,    1.85,
  2.33,    2.33,    2.33,    2.33,
  1.83,    1.83,    1.83,    1.83,
  2.31,    2.31,    2.31,    2.31,
  2.74,    2.74,    2.74,    2.74,
  2.88,    2.88,    2.88,    2.88,
  2.77,    2.77,    2.77,    2.77,
  2.84,    2.84,    2.84,    2.84,
  2.87,    2.87,    2.87,    2.87,
  2.58,    2.58,    2.58,    2.58,
  2.6,     2.6,     2.6,     2.6,
  2.86,    2.86,    2.86,    2.86,
  2.73,    2.73,    2.73,    2.73,
  2.53,    2.53,    2.53,    2.53,
  2.53,    2.53,    2.53,    2.53,
  2.42,    2.42,    2.42,    2.42,
  2.51,    2.51,    2.51,    2.51,
  2.41,    2.41,    2.41,    2.41,
  2.24,    2.24,    2.24,    2.24,
  1.91,    1.91,    1.91,    1.91,
  1.75,    1.75,    1.75,    1.75,
  1.7,     1.7,     1.7,     1.7,
  1.9,     1.9,     1.9,     1.9,
  1.56,    1.56,    1.56,    1.56,
  1.54,    1.54,    1.54,    1.54,
  1.93,    1.93,    1.93,    1.93,
  1.71,    1.71,    1.71,    1.71,
  1.51,    1.51,    1.51,    1.51,
  1.47,    1.47,    1.47,    1.47,
  2.03,    2.03,    2.03,    2.03,
  1.82,    1.82,    1.82,    1.82,
  1.59,    1.59,    1.59,    1.59,
  2.7,     2.7,     2.7,     2.7,
  2.24,    2.24,    2.24,    2.24,
  2.39,    2.39,    2.39,    2.39,
  2.53,    2.53,    2.53,    2.53,
  2.49,    2.49,    2.49,    2.49,
  2.3,     2.3,     2.3,     2.3,
  2.66,    2.66,    2.66,    2.66,
  3.06,    3.06,    3.06,    3.06,
  2.25,    2.25,    2.25,    2.25,
  1.92,    1.92,    1.92,    1.92,
  2.06,    2.06,    2.06,    2.06,
  2.14,    2.14,    2.14,    2.14,
  2.29,    2.29,    2.29,    2.29,
  2.76,    2.76,    2.76,    2.76,
  2.73,    2.73,    2.73,    2.73,
  2.68,    2.68,    2.68,    2.68,
  3.04,    3.04,    3.04,    3.04,
  4.07,    4.07,    4.07,    4.07,
  3.01,    3.01,    3.01,    3.01,
  1.79,    1.79,    1.79,    1.79,
  2.1,     2.1,     2.1,     2.1,
  2.53,    2.53,    2.53,    2.53,
  2.71,    2.71,    2.71,    2.71,
  2.78,    2.78,    2.78,    2.78,
  2.76,    2.76,    2.76,    2.76,
  3.18,    3.18,    3.18,    3.18,
  3,       3,       3,       3,
  3.33,    3.33,    3.33,    3.33,
  3.86,    3.86,    3.86,    3.86,
  3.07,    3.07,    3.07,    3.07,
  2.91,    2.91,    2.91,    2.91,
  3.05,    3.05,    3.05,    3.05,
  3.59,    3.59,    3.59,    3.59,
  3.76,    3.76,    3.76,    3.76,
  3.44,    3.44,    3.44,    3.44,
  3.73,    3.73,    3.73,    3.73,
  4.03,    4.03,    4.03,    4.03,
  3.86,    3.86,    3.86,    3.86,
  3.91,    3.91,    3.91,    3.91,
  3.98,    3.98,    3.98,    3.98,
  4.08,    4.08,    4.08,    4.08,
  3.53,    3.53,    3.53,    3.53,
  4.66,    4.66,    4.66,    4.66,
  4.44,    4.44,    4.44,    4.44,
  4.46,    4.46,    4.46,    4.46,
  4.64,    4.64,    4.64,    4.64,
  4.4,     4.4,     4.4,     4.4,
  5.22,    5.22,    5.22,    5.22,
  3.77,    3.77,    3.77,    3.77,
  5.37,    5.37,    5.37,    5.37,
  5.04,    5.04,    5.04,    5.04,
  5.37,    5.37,    5.37,    5.37,
  3.51,    3.51,    3.51,    3.51,
  3.39,    3.39,    3.39,    3.39,
  4.62,    4.62,    4.62,    4.62,
  3.2,     3.2,     3.2,     3.2,
  4.3,     4.3,     4.3,     4.3,
  4.52,    4.52,    4.52,    4.52,
  3.18,    3.18,    3.18,    3.18,
  3.62,    3.62,    3.62,    3.62,
  4,       4,       4,       4,
  4.22,    4.22,    4.22,    4.22,
  3.91,    3.91,    3.91,    3.91,
  3.48,    3.48,    3.48,    3.48,
  3.18,    3.18,    3.18,    3.18,
  2.18,    2.18,    2.18,    2.18,
  1.8,     1.8,     1.8,     1.8,
  0.75,    0.75,    0.75,    0.75,
  0.67,    0.67,    0.67,    0.67,
  1.88,    1.88,    1.88,    1.88,
  1.96,    1.96,    1.96,    1.96,
  1.99,    1.99,    1.99,    1.99,
  2.09,    2.09,    2.09,    2.09,
  2.11,    2.11,    2.11,    2.11,
  2.09,    2.09,    2.09,    2.09,
  2.29,    2.29,    2.29,    2.29,
  2.12,    2.12,    2.12,    2.12,
  2.25,    2.25,    2.25,    2.25,
  1.91,    1.91,    1.91,    1.91,
  2.21,    2.21,    2.21,    2.21,
  2.11,    2.11,    2.11,    2.11,
  2.14,    2.14,    2.14,    2.14,
  2.13,    2.13,    2.13,    2.13,
  2.19,    2.19,    2.19,    2.19,
  2.52,    2.52,    2.52,    2.52,
  2.26,    2.26,    2.26,    2.26,
  1.88,    1.88,    1.88,    1.88,
  1.83,    1.83,    1.83,    1.83,
  2.04,    2.04,    2.04,    2.04,
  1.99,    1.99,    1.99,    1.99,
  2.08,    2.08,    2.08,    2.08,
  2.48,    2.48,    2.48,    2.48,
  2.35,    2.35,    2.35,    2.35,
  2.21,    2.21,    2.21,    2.21,
  2.42,    2.42,    2.42,    2.42,
  2.24,    2.24,    2.24,    2.24,
  3.38,    3.38,    3.38,    3.38,
  2.66,    2.66,    2.66,    2.66,
  2.81,    2.81,    2.81,    2.81,
  2.43,    2.43,    2.43,    2.43,
  2.26,    2.26,    2.26,    2.26,
  2.63,    2.63,    2.63,    2.63,
  3.41,    3.41,    3.41,    3.41,
  3.79,    3.79,    3.79,    3.79,
  3.01,    3.01,    3.01,    3.01,
  3.28,    3.28,    3.28,    3.28,
  3.87,    3.87,    3.87,    3.87,
  3.58,    3.58,    3.58,    3.58,
  3.17,    3.17,    3.17,    3.17,
  2.64,    2.64,    2.64,    2.64,
  2.83,    2.83,    2.83,    2.83,
  2.36,    2.36,    2.36,    2.36,
  2.24,    2.24,    2.24,    2.24,
  2.28,    2.28,    2.28,    2.28,
  2.64,    2.64,    2.64,    2.64,
  2.21,    2.21,    2.21,    2.21,
  2.21,    2.21,    2.21,    2.21,
  2.32,    2.32,    2.32,    2.32,
  1.8,     1.8,     1.8,     1.8,
  1.84,    1.84,    1.84,    1.84,
  2.34,    2.34,    2.34,    2.34,
  2.41,    2.41,    2.41,    2.41,
  2.37,    2.37,    2.37,    2.37,
  2.4,     2.4,     2.4,     2.4,
  2.49,    2.49,    2.49,    2.49,
  2.34,    2.34,    2.34,    2.34,
  2.4,     2.4,     2.4,     2.4,
  2.79,    2.79,    2.79,    2.79,
  3.12,    3.12,    3.12,    3.12,
  2.4,     2.4,     2.4,     2.4,
  2.36,    2.36,    2.36,    2.36,
  1.9,     1.9,     1.9,     1.9,
  1.92,    1.92,    1.92,    1.92,
  1.5,     1.5,     1.5,     1.5,
  1.55,    1.55,    1.55,    1.55,
  1.42,    1.42,    1.42,    1.42,
  1.38,    1.38,    1.38,    1.38,
  1.39,    1.39,    1.39,    1.39,
  1.57,    1.57,    1.57,    1.57,
  1.56,    1.56,    1.56,    1.56,
  1.89,    1.89,    1.89,    1.89,
  2.18,    2.18,    2.18,    2.18,
  2.1,     2.1,     2.1,     2.1,
  2.13,    2.13,    2.13,    2.13,
  2.07,    2.07,    2.07,    2.07,
  2.06,    2.06,    2.06,    2.06,
  2.61,    2.61,    2.61,    2.61,
  2.51,    2.51,    2.51,    2.51,
  2.62,    2.62,    2.62,    2.62,
  3.07,    3.07,    3.07,    3.07,
  2.61,    2.61,    2.61,    2.61,
  3,       3,       3,       3,
  3.2,     3.2,     3.2,     3.2,
  2.93,    2.93,    2.93,    2.93,
  2.36,    2.36,    2.36,    2.36,
  2.85,    2.85,    2.85,    2.85,
  3.13,    3.13,    3.13,    3.13,
  3.38,    3.38,    3.38,    3.38,
  2.81,    2.81,    2.81,    2.81,
  2.66,    2.66,    2.66,    2.66,
  2.49,    2.49,    2.49,    2.49,
  2.35,    2.35,    2.35,    2.35,
  2.92,    2.92,    2.92,    2.92,
  2.85,    2.85,    2.85,    2.85,
  2.85,    2.85,    2.85,    2.85,
  2.85,    2.85,    2.85,    2.85,
  2.96,    2.96,    2.96,    2.96,
  2.46,    2.46,    2.46,    2.46,
  2.5,     2.5,     2.5,     2.5,
  2.94,    2.94,    2.94,    2.94,
  2.71,    2.71,    2.71,    2.71,
  2.52,    2.52,    2.52,    2.52,
  2.57,    2.57,    2.57,    2.57,
  2.44,    2.44,    2.44,    2.44,
  2.27,    2.27,    2.27,    2.27,
  2.34,    2.34,    2.34,    2.34,
  2.09,    2.09,    2.09,    2.09,
  1.85,    1.85,    1.85,    1.85,
  1.83,    1.83,    1.83,    1.83,
  1.93,    1.93,    1.93,    1.93,
  2.03,    2.03,    2.03,    2.03,
  2.12,    2.12,    2.12,    2.12,
  2.41,    2.41,    2.41,    2.41,
  2.21,    2.21,    2.21,    2.21,
  2.18,    2.18,    2.18,    2.18,
  2.48,    2.48,    2.48,    2.48,
  2.39,    2.39,    2.39,    2.39,
  2.59,    2.59,    2.59,    2.59,
  2.9,     2.9,     2.9,     2.9,
  2.73,    2.73,    2.73,    2.73,
  2.99,    2.99,    2.99,    2.99,
  3.54,    3.54,    3.54,    3.54,
  2.97,    2.97,    2.97,    2.97,
  3.26,    3.26,    3.26,    3.26,
  3.1,     3.1,     3.1,     3.1,
  3.93,    3.93,    3.93,    3.93,
  4.45,    4.45,    4.45,    4.45,
  3.19,    3.19,    3.19,    3.19,
  3.22,    3.22,    3.22,    3.22,
  3.34,    3.34,    3.34,    3.34,
  2.98,    2.98,    2.98,    2.98,
  3.32,    3.32,    3.32,    3.32,
  3.2,     3.2,     3.2,     3.2,
  2.22,    2.22,    2.22,    2.22,
  1.15,    1.15,    1.15,    1.15,
  1.28,    1.28,    1.28,    1.28,
  1.51,    1.51,    1.51,    1.51,
  1.52,    1.52,    1.52,    1.52,
  1.43,    1.43,    1.43,    1.43,
  1.55,    1.55,    1.55,    1.55,
  2.23,    2.23,    2.23,    2.23,
  2.14,    2.14,    2.14,    2.14,
  2.03,    2.03,    2.03,    2.03,
  1.85,    1.85,    1.85,    1.85,
  1.93,    1.93,    1.93,    1.93,
  1.85,    1.85,    1.85,    1.85,
  1.72,    1.72,    1.72,    1.72,
  2.32,    2.32,    2.32,    2.32,
  2.48,    2.48,    2.48,    2.48,
  2.03,    2.03,    2.03,    2.03,
  1.96,    1.96,    1.96,    1.96,
  2.26,    2.26,    2.26,    2.26,
  2.04,    2.04,    2.04,    2.04,
  2.19,    2.19,    2.19,    2.19,
  1.77,    1.77,    1.77,    1.77,
  1.61,    1.61,    1.61,    1.61,
  1.58,    1.58,    1.58,    1.58,
  1.17,    1.17,    1.17,    1.17,
  1.08,    1.08,    1.08,    1.08,
  0.94,    0.94,    0.94,    0.94,
  1.19,    1.19,    1.19,    1.19,
  1.14,    1.14,    1.14,    1.14,
  0.65,    0.65,    0.65,    0.65,
  0.29,    0.29,    0.29,    0.29,
  0.17,    0.17,    0.17,    0.17,
  0.99,    0.99,    0.99,    0.99,
  1.12,    1.12,    1.12,    1.12,
  1,       1,       1,       1,
  1.03,    1.03,    1.03,    1.03,
  1.25,    1.25,    1.25,    1.25,
  0.88,    0.88,    0.88,    0.88,
  1.42,    1.42,    1.42,    1.42,
  1.61,    1.61,    1.61,    1.61,
  0.25,    0.25,    0.25,    0.25,
  0.96,    0.96,    0.96,    0.96,
  1.68,    1.68,    1.68,    1.68,
  1.48,    1.48,    1.48,    1.48,
  1.45,    1.45,    1.45,    1.45,
  1.67,    1.67,    1.67,    1.67,
  1.72,    1.72,    1.72,    1.72,
  0.79,    0.79,    0.79,    0.79,
  0.83,    0.83,    0.83,    0.83,
  0.68,    0.68,    0.68,    0.68,
  1.24,    1.24,    1.24,    1.24,
  1.12,    1.12,    1.12,    1.12,
  1.9,     1.9,     1.9,     1.9,
  1.43,    1.43,    1.43,    1.43,
  1.73,    1.73,    1.73,    1.73,
  2.03,    2.03,    2.03,    2.03,
  2.05,    2.05,    2.05,    2.05,
  2.09,    2.09,    2.09,    2.09,
  1.88,    1.88,    1.88,    1.88,
  1.64,    1.64,    1.64,    1.64,
  1.77,    1.77,    1.77,    1.77,
  1.87,    1.87,    1.87,    1.87,
  1.9,     1.9,     1.9,     1.9,
  1.67,    1.67,    1.67,    1.67,
  1.87,    1.87,    1.87,    1.87,
  1.91,    1.91,    1.91,    1.91,
  1.81,    1.81,    1.81,    1.81,
  1.96,    1.96,    1.96,    1.96,
  2.2,     2.2,     2.2,     2.2,
  2.11,    2.11,    2.11,    2.11,
  2.04,    2.04,    2.04,    2.04,
  1.84,    1.84,    1.84,    1.84,
  1.77,    1.77,    1.77,    1.77,
  1.99,    1.99,    1.99,    1.99,
  2.13,    2.13,    2.13,    2.13,
  1.83,    1.83,    1.83,    1.83,
  1.9,     1.9,     1.9,     1.9,
  2.27,    2.27,    2.27,    2.27,
  1.99,    1.99,    1.99,    1.99,
  1.6,     1.6,     1.6,     1.6,
  1.3,     1.3,     1.3,     1.3,
  1.29,    1.29,    1.29,    1.29,
  2.04,    2.04,    2.04,    2.04,
  2.55,    2.55,    2.55,    2.55,
  2.54,    2.54,    2.54,    2.54,
  2.31,    2.31,    2.31,    2.31,
  2.03,    2.03,    2.03,    2.03,
  1.89,    1.89,    1.89,    1.89,
  2.11,    2.11,    2.11,    2.11,
  2.82,    2.82,    2.82,    2.82,
  1.95,    1.95,    1.95,    1.95,
  2.26,    2.26,    2.26,    2.26,
  2.38,    2.38,    2.38,    2.38,
  2.43,    2.43,    2.43,    2.43,
  2.51,    2.51,    2.51,    2.51,
  2.04,    2.04,    2.04,    2.04,
  1.63,    1.63,    1.63,    1.63,
  2.37,    2.37,    2.37,    2.37,
  1.69,    1.69,    1.69,    1.69,
  1,       1,       1,       1,
  1.2,     1.2,     1.2,     1.2,
  1.56,    1.56,    1.56,    1.56,
  1.93,    1.93,    1.93,    1.93,
  1.83,    1.83,    1.83,    1.83,
  2.1,     2.1,     2.1,     2.1,
  2.05,    2.05,    2.05,    2.05,
  2.19,    2.19,    2.19,    2.19,
  2.23,    2.23,    2.23,    2.23,
  2.1,     2.1,     2.1,     2.1,
  2.02,    2.02,    2.02,    2.02,
  2.08,    2.08,    2.08,    2.08,
  2.05,    2.05,    2.05,    2.05,
  1.97,    1.97,    1.97,    1.97,
  2.08,    2.08,    2.08,    2.08,
  1.26,    1.26,    1.26,    1.26,
  1.87,    1.87,    1.87,    1.87,
  1.9,     1.9,     1.9,     1.9,
  1.85,    1.85,    1.85,    1.85,
  1.67,    1.67,    1.67,    1.67,
  1.79,    1.79,    1.79,    1.79,
  1.81,    1.81,    1.81,    1.81,
  1.69,    1.69,    1.69,    1.69,
  2.16,    2.16,    2.16,    2.16,
  2.07,    2.07,    2.07,    2.07,
  2.09,    2.09,    2.09,    2.09,
  1.3,     1.3,     1.3,     1.3,
  1.36,    1.36,    1.36,    1.36,
  0.56,    0.56,    0.56,    0.56,
  1.8,     1.8,     1.8,     1.8,
  2.12,    2.12,    2.12,    2.12,
  1.91,    1.91,    1.91,    1.91,
  2.13,    2.13,    2.13,    2.13,
  2.52,    2.52,    2.52,    2.52,
  1.97,    1.97,    1.97,    1.97,
  2.35,    2.35,    2.35,    2.35,
  2.47,    2.47,    2.47,    2.47,
  2.61,    2.61,    2.61,    2.61,
  2.8,     2.8,     2.8,     2.8,
  2.74,    2.74,    2.74,    2.74,
  3.37,    3.37,    3.37,    3.37,
  3.43,    3.43,    3.43,    3.43,
  3.55,    3.55,    3.55,    3.55,
  3.1,     3.1,     3.1,     3.1,
  3.07,    3.07,    3.07,    3.07,
  2.68,    2.68,    2.68,    2.68,
  2.56,    2.56,    2.56,    2.56,
  2.53,    2.53,    2.53,    2.53,
  2.16,    2.16,    2.16,    2.16,
  2.13,    2.13,    2.13,    2.13,
  1.36,    1.36,    1.36,    1.36,
  1.75,    1.75,    1.75,    1.75,
  1.84,    1.84,    1.84,    1.84,
  1.93,    1.93,    1.93,    1.93,
  1.82,    1.82,    1.82,    1.82,
  2.37,    2.37,    2.37,    2.37,
  1.68,    1.68,    1.68,    1.68,
  1.6,     1.6,     1.6,     1.6,
  1.63,    1.63,    1.63,    1.63,
  1.73,    1.73,    1.73,    1.73,
  1.75,    1.75,    1.75,    1.75,
  1.35,    1.35,    1.35,    1.35,
  1.12,    1.12,    1.12,    1.12,
  1.58,    1.58,    1.58,    1.58,
  1.03,    1.03,    1.03,    1.03,
  1.35,    1.35,    1.35,    1.35,
  1.6,     1.6,     1.6,     1.6,
  1.52,    1.52,    1.52,    1.52,
  1.2,     1.2,     1.2,     1.2,
  1.63,    1.63,    1.63,    1.63,
  1.26,    1.26,    1.26,    1.26,
  1.44,    1.44,    1.44,    1.44,
  1.12,    1.12,    1.12,    1.12,
  0.47,    0.47,    0.47,    0.47,
  0.86,    0.86,    0.86,    0.86,
  0.28,    0.28,    0.28,    0.28,
  0.6,     0.6,     0.6,     0.6,
  0.84,    0.84,    0.84,    0.84,
  1.26,    1.26,    1.26,    1.26,
  0.96,    0.96,    0.96,    0.96,
  1.34,    1.34,    1.34,    1.34,
  1.54,    1.54,    1.54,    1.54,
  1.64,    1.64,    1.64,    1.64,
  1.81,    1.81,    1.81,    1.81,
  1.71,    1.71,    1.71,    1.71,
  1.56,    1.56,    1.56,    1.56,
  2.08,    2.08,    2.08,    2.08,
  1.89,    1.89,    1.89,    1.89,
  1.64,    1.64,    1.64,    1.64,
  1.39,    1.39,    1.39,    1.39,
  1.2,     1.2,     1.2,     1.2,
  1.85,    1.85,    1.85,    1.85,
  1.85,    1.85,    1.85,    1.85,
  2.12,    2.12,    2.12,    2.12,
  1.55,    1.55,    1.55,    1.55,
  1.23,    1.23,    1.23,    1.23,
  1.76,    1.76,    1.76,    1.76,
  1.49,    1.49,    1.49,    1.49,
  1.56,    1.56,    1.56,    1.56,
  1.83,    1.83,    1.83,    1.83,
  1.15,    1.15,    1.15,    1.15,
  1.41,    1.41,    1.41,    1.41,
  1.4,     1.4,     1.4,     1.4,
  2,       2,       2,       2,
  2.07,    2.07,    2.07,    2.07,
  1.88,    1.88,    1.88,    1.88,
  1.84,    1.84,    1.84,    1.84,
  1.81,    1.81,    1.81,    1.81,
  2.13,    2.13,    2.13,    2.13,
  2.43,    2.43,    2.43,    2.43,
  2.35,    2.35,    2.35,    2.35,
  2.16,    2.16,    2.16,    2.16,
  2.02,    2.02,    2.02,    2.02,
  2.04,    2.04,    2.04,    2.04,
  2.24,    2.24,    2.24,    2.24,
  2.02,    2.02,    2.02,    2.02,
  1.59,    1.59,    1.59,    1.59,
  1.55,    1.55,    1.55,    1.55,
  1.64,    1.64,    1.64,    1.64,
  2.02,    2.02,    2.02,    2.02,
  2.03,    2.03,    2.03,    2.03,
  1.82,    1.82,    1.82,    1.82,
  1.36,    1.36,    1.36,    1.36,
  1.41,    1.41,    1.41,    1.41,
  1.3,     1.3,     1.3,     1.3,
  1.43,    1.43,    1.43,    1.43,
  2.26,    2.26,    2.26,    2.26,
  2.73,    2.73,    2.73,    2.73,
  2.46,    2.46,    2.46,    2.46,
  2.59,    2.59,    2.59,    2.59,
  1.89,    1.89,    1.89,    1.89,
  3.02,    3.02,    3.02,    3.02,
  3.55,    3.55,    3.55,    3.55,
  3.48,    3.48,    3.48,    3.48,
  3.91,    3.91,    3.91,    3.91,
  4.62,    4.62,    4.62,    4.62,
  4.2,     4.2,     4.2,     4.2,
  5.18,    5.18,    5.18,    5.18,
  4.96,    4.96,    4.96,    4.96,
  4.69,    4.69,    4.69,    4.69,
  4.93,    4.93,    4.93,    4.93,
  4.93,    4.93,    4.93,    4.93,
  4.55,    4.55,    4.55,    4.55,
  4.23,    4.23,    4.23,    4.23,
  3.52,    3.52,    3.52,    3.52,
  2.82,    2.82,    2.82,    2.82,
  2.12,    2.12,    2.12,    2.12,
  2.26,    2.26,    2.26,    2.26,
  2.12,    2.12,    2.12,    2.12,
  2.08,    2.08,    2.08,    2.08,
  2.23,    2.23,    2.23,    2.23,
  2.21,    2.21,    2.21,    2.21,
  2.21,    2.21,    2.21,    2.21,
  2.23,    2.23,    2.23,    2.23,
  2.51,    2.51,    2.51,    2.51,
  2.53,    2.53,    2.53,    2.53,
  2.52,    2.52,    2.52,    2.52,
  2.41,    2.41,    2.41,    2.41,
  2,       2,       2,       2,
  2.02,    2.02,    2.02,    2.02,
  1.86,    1.86,    1.86,    1.86,
  1.75,    1.75,    1.75,    1.75,
  1.87,    1.87,    1.87,    1.87,
  2.09,    2.09,    2.09,    2.09,
  2.46,    2.46,    2.46,    2.46,
  2.74,    2.74,    2.74,    2.74,
  2.72,    2.72,    2.72,    2.72,
  2.97,    2.97,    2.97,    2.97,
  3.11,    3.11,    3.11,    3.11,
  3.11,    3.11,    3.11,    3.11,
  3.26,    3.26,    3.26,    3.26,
  2.84,    2.84,    2.84,    2.84,
  2.18,    2.18,    2.18,    2.18,
  2.66,    2.66,    2.66,    2.66,
  2.26,    2.26,    2.26,    2.26,
  1.93,    1.93,    1.93,    1.93,
  2.16,    2.16,    2.16,    2.16,
  2.4,     2.4,     2.4,     2.4,
  2.05,    2.05,    2.05,    2.05,
  2.6,     2.6,     2.6,     2.6,
  2.58,    2.58,    2.58,    2.58,
  2.13,    2.13,    2.13,    2.13,
  1.99,    1.99,    1.99,    1.99,
  2.71,    2.71,    2.71,    2.71,
  3.5,     3.5,     3.5,     3.5,
  3.71,    3.71,    3.71,    3.71,
  3.54,    3.54,    3.54,    3.54,
  4.13,    4.13,    4.13,    4.13,
  3.75,    3.75,    3.75,    3.75,
  3.98,    3.98,    3.98,    3.98,
  3.86,    3.86,    3.86,    3.86,
  3.43,    3.43,    3.43,    3.43,
  2.96,    2.96,    2.96,    2.96,
  2.68,    2.68,    2.68,    2.68,
  2.14,    2.14,    2.14,    2.14,
  2.3,     2.3,     2.3,     2.3,
  2.12,    2.12,    2.12,    2.12,
  2.14,    2.14,    2.14,    2.14,
  1.75,    1.75,    1.75,    1.75,
  1.82,    1.82,    1.82,    1.82,
  2.04,    2.04,    2.04,    2.04,
  2.19,    2.19,    2.19,    2.19,
  2.18,    2.18,    2.18,    2.18,
  2.33,    2.33,    2.33,    2.33,
  2.37,    2.37,    2.37,    2.37,
  2.3,     2.3,     2.3,     2.3,
  2.43,    2.43,    2.43,    2.43,
  2.38,    2.38,    2.38,    2.38,
  2.4,     2.4,     2.4,     2.4,
  2.21,    2.21,    2.21,    2.21,
  2.32,    2.32,    2.32,    2.32,
  2.28,    2.28,    2.28,    2.28,
  2.34,    2.34,    2.34,    2.34,
  2.67,    2.67,    2.67,    2.67,
  3.01,    3.01,    3.01,    3.01,
  2.85,    2.85,    2.85,    2.85,
  2.63,    2.63,    2.63,    2.63,
  2.66,    2.66,    2.66,    2.66,
  2.54,    2.54,    2.54,    2.54,
  2.47,    2.47,    2.47,    2.47,
  2.54,    2.54,    2.54,    2.54,
  2.9,     2.9,     2.9,     2.9,
  3.02,    3.02,    3.02,    3.02,
  4.54,    4.54,    4.54,    4.54,
  4.36,    4.36,    4.36,    4.36,
  4.65,    4.65,    4.65,    4.65,
  4.79,    4.79,    4.79,    4.79,
  4.83,    4.83,    4.83,    4.83,
  5.23,    5.23,    5.23,    5.23,
  5.14,    5.14,    5.14,    5.14,
  4.59,    4.59,    4.59,    4.59,
  4.81,    4.81,    4.81,    4.81,
  4.6,     4.6,     4.6,     4.6,
  4.59,    4.59,    4.59,    4.59,
  4.86,    4.86,    4.86,    4.86,
  4.22,    4.22,    4.22,    4.22,
  4.34,    4.34,    4.34,    4.34,
  4.21,    4.21,    4.21,    4.21,
  3.76,    3.76,    3.76,    3.76,
  3.41,    3.41,    3.41,    3.41,
  3.61,    3.61,    3.61,    3.61,
  3.81,    3.81,    3.81,    3.81,
  3.1,     3.1,     3.1,     3.1,
  2.66,    2.66,    2.66,    2.66,
  2.07,    2.07,    2.07,    2.07,
  2.05,    2.05,    2.05,    2.05,
  2.36,    2.36,    2.36,    2.36,
  2.23,    2.23,    2.23,    2.23,
  1.81,    1.81,    1.81,    1.81,
  1.79,    1.79,    1.79,    1.79,
  1.8,     1.8,     1.8,     1.8,
  2.51,    2.51,    2.51,    2.51,
  2.47,    2.47,    2.47,    2.47,
  2.39,    2.39,    2.39,    2.39,
  2.45,    2.45,    2.45,    2.45,
  2.55,    2.55,    2.55,    2.55,
  1.72,    1.72,    1.72,    1.72,
  1.86,    1.86,    1.86,    1.86,
  1.67,    1.67,    1.67,    1.67,
  1.69,    1.69,    1.69,    1.69,
  1.79,    1.79,    1.79,    1.79,
  1.97,    1.97,    1.97,    1.97,
  2.09,    2.09,    2.09,    2.09,
  2.36,    2.36,    2.36,    2.36,
  1.96,    1.96,    1.96,    1.96,
  1.77,    1.77,    1.77,    1.77,
  1.98,    1.98,    1.98,    1.98,
  1.76,    1.76,    1.76,    1.76,
  1.91,    1.91,    1.91,    1.91,
  2.34,    2.34,    2.34,    2.34,
  2.93,    2.93,    2.93,    2.93,
  3.62,    3.62,    3.62,    3.62,
  4.22,    4.22,    4.22,    4.22,
  4.52,    4.52,    4.52,    4.52,
  4.45,    4.45,    4.45,    4.45,
  4.54,    4.54,    4.54,    4.54,
  6.04,    6.04,    6.04,    6.04,
  5.81,    5.81,    5.81,    5.81,
  6.16,    6.16,    6.16,    6.16,
  5.53,    5.53,    5.53,    5.53,
  5.49,    5.49,    5.49,    5.49,
  6.3,     6.3,     6.3,     6.3,
  5.86,    5.86,    5.86,    5.86,
  5.85,    5.85,    5.85,    5.85,
  4.9,     4.9,     4.9,     4.9,
  5.59,    5.59,    5.59,    5.59,
  4.93,    4.93,    4.93,    4.93,
  5.39,    5.39,    5.39,    5.39,
  4.56,    4.56,    4.56,    4.56,
  4.09,    4.09,    4.09,    4.09,
  4.11,    4.11,    4.11,    4.11,
  3.95,    3.95,    3.95,    3.95,
  4.71,    4.71,    4.71,    4.71,
  3.09,    3.09,    3.09,    3.09,
  2.92,    2.92,    2.92,    2.92,
  2.59,    2.59,    2.59,    2.59,
  1.84,    1.84,    1.84,    1.84,
  1.84,    1.84,    1.84,    1.84,
  1.82,    1.82,    1.82,    1.82,
  2.4,     2.4,     2.4,     2.4,
  2.94,    2.94,    2.94,    2.94,
  2.42,    2.42,    2.42,    2.42,
  2.54,    2.54,    2.54,    2.54,
  2.32,    2.32,    2.32,    2.32,
  1.81,    1.81,    1.81,    1.81,
  1.73,    1.73,    1.73,    1.73,
  1.56,    1.56,    1.56,    1.56,
  1.68,    1.68,    1.68,    1.68,
  1.76,    1.76,    1.76,    1.76,
  1.73,    1.73,    1.73,    1.73,
  2.14,    2.14,    2.14,    2.14,
  1.8,     1.8,     1.8,     1.8,
  1.75,    1.75,    1.75,    1.75,
  1.98,    1.98,    1.98,    1.98,
  1.87,    1.87,    1.87,    1.87,
  1.5,     1.5,     1.5,     1.5,
  1.46,    1.46,    1.46,    1.46,
  1.94,    1.94,    1.94,    1.94,
  2.7,     2.7,     2.7,     2.7,
  3.05,    3.05,    3.05,    3.05,
  2.89,    2.89,    2.89,    2.89,
  2.95,    2.95,    2.95,    2.95,
  3.03,    3.03,    3.03,    3.03,
  2.71,    2.71,    2.71,    2.71,
  2.82,    2.82,    2.82,    2.82,
  2.66,    2.66,    2.66,    2.66,
  2.99,    2.99,    2.99,    2.99,
  2.95,    2.95,    2.95,    2.95,
  3.02,    3.02,    3.02,    3.02,
  2.84,    2.84,    2.84,    2.84,
  2.01,    2.01,    2.01,    2.01,
  3.32,    3.32,    3.32,    3.32,
  2.1,     2.1,     2.1,     2.1,
  2.24,    2.24,    2.24,    2.24,
  2.2,     2.2,     2.2,     2.2,
  2.07,    2.07,    2.07,    2.07,
  1.98,    1.98,    1.98,    1.98,
  1.72,    1.72,    1.72,    1.72,
  1.57,    1.57,    1.57,    1.57,
  1.77,    1.77,    1.77,    1.77,
  1.81,    1.81,    1.81,    1.81,
  1.31,    1.31,    1.31,    1.31,
  1.49,    1.49,    1.49,    1.49,
  1.47,    1.47,    1.47,    1.47,
  1.81,    1.81,    1.81,    1.81,
  2.24,    2.24,    2.24,    2.24,
  2.04,    2.04,    2.04,    2.04,
  2.03,    2.03,    2.03,    2.03,
  1.94,    1.94,    1.94,    1.94,
  1.27,    1.27,    1.27,    1.27,
  2.46,    2.46,    2.46,    2.46,
  2.25,    2.25,    2.25,    2.25,
  2.44,    2.44,    2.44,    2.44,
  2.69,    2.69,    2.69,    2.69,
  2.56,    2.56,    2.56,    2.56,
  2.19,    2.19,    2.19,    2.19,
  2.33,    2.33,    2.33,    2.33,
  2.47,    2.47,    2.47,    2.47,
  2.51,    2.51,    2.51,    2.51,
  2.08,    2.08,    2.08,    2.08,
  1.64,    1.64,    1.64,    1.64,
  2.12,    2.12,    2.12,    2.12,
  2.36,    2.36,    2.36,    2.36,
  2.52,    2.52,    2.52,    2.52,
  2.29,    2.29,    2.29,    2.29,
  2.17,    2.17,    2.17,    2.17,
  2.09,    2.09,    2.09,    2.09,
  3.45,    3.45,    3.45,    3.45,
  3.1,     3.1,     3.1,     3.1,
  2.7,     2.7,     2.7,     2.7,
  2.66,    2.66,    2.66,    2.66,
  2.86,    2.86,    2.86,    2.86,
  2.62,    2.62,    2.62,    2.62,
  3.58,    3.58,    3.58,    3.58,
  3.35,    3.35,    3.35,    3.35,
  3.2,     3.2,     3.2,     3.2,
  3.09,    3.09,    3.09,    3.09,
  2.86,    2.86,    2.86,    2.86,
  2.93,    2.93,    2.93,    2.93,
  3.69,    3.69,    3.69,    3.69,
  3.66,    3.66,    3.66,    3.66,
  2.63,    2.63,    2.63,    2.63,
  2.44,    2.44,    2.44,    2.44,
  1.79,    1.79,    1.79,    1.79,
  1.89,    1.89,    1.89,    1.89,
  2.22,    2.22,    2.22,    2.22,
  2.29,    2.29,    2.29,    2.29,
  2.12,    2.12,    2.12,    2.12,
  2.17,    2.17,    2.17,    2.17,
  2.33,    2.33,    2.33,    2.33,
  2.51,    2.51,    2.51,    2.51,
  2.53,    2.53,    2.53,    2.53,
  2.81,    2.81,    2.81,    2.81,
  2.88,    2.88,    2.88,    2.88,
  2.69,    2.69,    2.69,    2.69,
  2.77,    2.77,    2.77,    2.77,
  2.73,    2.73,    2.73,    2.73,
  2.44,    2.44,    2.44,    2.44,
  2.47,    2.47,    2.47,    2.47,
  2.39,    2.39,    2.39,    2.39,
  2.47,    2.47,    2.47,    2.47,
  2.66,    2.66,    2.66,    2.66,
  2.85,    2.85,    2.85,    2.85,
  3.1,     3.1,     3.1,     3.1,
  3.1,     3.1,     3.1,     3.1,
  2.99,    2.99,    2.99,    2.99,
  2.96,    2.96,    2.96,    2.96,
  2.99,    2.99,    2.99,    2.99,
  3.25,    3.25,    3.25,    3.25,
  3.36,    3.36,    3.36,    3.36,
  2.85,    2.85,    2.85,    2.85,
  3.09,    3.09,    3.09,    3.09,
  3.28,    3.28,    3.28,    3.28,
  3.85,    3.85,    3.85,    3.85,
  4.24,    4.24,    4.24,    4.24,
  4.59,    4.59,    4.59,    4.59,
  5.15,    5.15,    5.15,    5.15,
  4.76,    4.76,    4.76,    4.76,
  5.5,     5.5,     5.5,     5.5,
  5.39,    5.39,    5.39,    5.39,
  5.15,    5.15,    5.15,    5.15,
  4.9,     4.9,     4.9,     4.9,
  4.99,    4.99,    4.99,    4.99,
  4.61,    4.61,    4.61,    4.61,
  4.52,    4.52,    4.52,    4.52,
  4.38,    4.38,    4.38,    4.38,
  3.51,    3.51,    3.51,    3.51,
  3.64,    3.64,    3.64,    3.64,
  4.09,    4.09,    4.09,    4.09,
  3.23,    3.23,    3.23,    3.23,
  3.17,    3.17,    3.17,    3.17,
  3.44,    3.44,    3.44,    3.44,
  4.49,    4.49,    4.49,    4.49,
  4.62,    4.62,    4.62,    4.62,
  4.43,    4.43,    4.43,    4.43,
  4.71,    4.71,    4.71,    4.71,
  5.18,    5.18,    5.18,    5.18,
  5.03,    5.03,    5.03,    5.03,
  4.2,     4.2,     4.2,     4.2,
  3.37,    3.37,    3.37,    3.37,
  2.81,    2.81,    2.81,    2.81,
  2.76,    2.76,    2.76,    2.76,
  2.45,    2.45,    2.45,    2.45,
  1.82,    1.82,    1.82,    1.82,
  2.1,     2.1,     2.1,     2.1,
  1.68,    1.68,    1.68,    1.68,
  1.72,    1.72,    1.72,    1.72,
  2.01,    2.01,    2.01,    2.01,
  2.24,    2.24,    2.24,    2.24,
  2.26,    2.26,    2.26,    2.26,
  1.95,    1.95,    1.95,    1.95,
  1.91,    1.91,    1.91,    1.91,
  2.05,    2.05,    2.05,    2.05,
  2.28,    2.28,    2.28,    2.28,
  2.67,    2.67,    2.67,    2.67,
  2.86,    2.86,    2.86,    2.86,
  2.76,    2.76,    2.76,    2.76,
  2.63,    2.63,    2.63,    2.63,
  2.75,    2.75,    2.75,    2.75,
  2.78,    2.78,    2.78,    2.78,
  2.92,    2.92,    2.92,    2.92,
  3.58,    3.58,    3.58,    3.58,
  3.22,    3.22,    3.22,    3.22,
  3.88,    3.88,    3.88,    3.88,
  4.16,    4.16,    4.16,    4.16,
  3.8,     3.8,     3.8,     3.8,
  4.34,    4.34,    4.34,    4.34,
  5.39,    5.39,    5.39,    5.39,
  5.79,    5.79,    5.79,    5.79,
  6.6,     6.6,     6.6,     6.6,
  5.73,    5.73,    5.73,    5.73,
  6.43,    6.43,    6.43,    6.43,
  5.48,    5.48,    5.48,    5.48,
  6.32,    6.32,    6.32,    6.32,
  6.34,    6.34,    6.34,    6.34,
  6.61,    6.61,    6.61,    6.61,
  5.7,     5.7,     5.7,     5.7,
  5.72,    5.72,    5.72,    5.72,
  3.52,    3.52,    3.52,    3.52,
  3.52,    3.52,    3.52,    3.52,
  2.78,    2.78,    2.78,    2.78,
  2.19,    2.19,    2.19,    2.19,
  2.24,    2.24,    2.24,    2.24,
  2,       2,       2,       2,
  1.71,    1.71,    1.71,    1.71,
  2.16,    2.16,    2.16,    2.16,
  0.21,    0.21,    0.21,    0.21,
  2.24,    2.24,    2.24,    2.24,
  2.22,    2.22,    2.22,    2.22,
  2.94,    2.94,    2.94,    2.94,
  3.05,    3.05,    3.05,    3.05,
  2.74,    2.74,    2.74,    2.74,
  2.65,    2.65,    2.65,    2.65,
  2.47,    2.47,    2.47,    2.47,
  3.12,    3.12,    3.12,    3.12,
  2.86,    2.86,    2.86,    2.86,
  3,       3,       3,       3,
  2.81,    2.81,    2.81,    2.81,
  2.57,    2.57,    2.57,    2.57,
  3.15,    3.15,    3.15,    3.15,
  3.27,    3.27,    3.27,    3.27,
  2.59,    2.59,    2.59,    2.59,
  2.24,    2.24,    2.24,    2.24,
  1.75,    1.75,    1.75,    1.75,
  2.1,     2.1,     2.1,     2.1,
  1.79,    1.79,    1.79,    1.79,
  2.15,    2.15,    2.15,    2.15,
  2.29,    2.29,    2.29,    2.29,
  2.77,    2.77,    2.77,    2.77,
  2.71,    2.71,    2.71,    2.71,
  3.54,    3.54,    3.54,    3.54,
  3.32,    3.32,    3.32,    3.32,
  3.93,    3.93,    3.93,    3.93,
  3.96,    3.96,    3.96,    3.96,
  3.7,     3.7,     3.7,     3.7,
  3.77,    3.77,    3.77,    3.77,
  4.15,    4.15,    4.15,    4.15,
  4.3,     4.3,     4.3,     4.3,
  4.28,    4.28,    4.28,    4.28,
  4.28,    4.28,    4.28,    4.28,
  4.46,    4.46,    4.46,    4.46,
  3.76,    3.76,    3.76,    3.76,
  3.57,    3.57,    3.57,    3.57,
  3.33,    3.33,    3.33,    3.33,
  4.64,    4.64,    4.64,    4.64,
  3.56,    3.56,    3.56,    3.56,
  3.51,    3.51,    3.51,    3.51,
  2.79,    2.79,    2.79,    2.79,
  2.48,    2.48,    2.48,    2.48,
  2.6,     2.6,     2.6,     2.6,
  2.04,    2.04,    2.04,    2.04,
  1.8,     1.8,     1.8,     1.8,
  2.16,    2.16,    2.16,    2.16,
  2.22,    2.22,    2.22,    2.22,
  2.32,    2.32,    2.32,    2.32,
  2.34,    2.34,    2.34,    2.34,
  2.23,    2.23,    2.23,    2.23,
  2.28,    2.28,    2.28,    2.28,
  2.28,    2.28,    2.28,    2.28,
  2.17,    2.17,    2.17,    2.17,
  2.26,    2.26,    2.26,    2.26,
  2.22,    2.22,    2.22,    2.22,
  2.21,    2.21,    2.21,    2.21,
  2.31,    2.31,    2.31,    2.31,
  2.2,     2.2,     2.2,     2.2,
  2.06,    2.06,    2.06,    2.06,
  2.08,    2.08,    2.08,    2.08,
  1.98,    1.98,    1.98,    1.98,
  1.92,    1.92,    1.92,    1.92,
  1.96,    1.96,    1.96,    1.96,
  2.08,    2.08,    2.08,    2.08,
  2.17,    2.17,    2.17,    2.17,
  2.11,    2.11,    2.11,    2.11,
  2.31,    2.31,    2.31,    2.31,
  2.51,    2.51,    2.51,    2.51,
  2.53,    2.53,    2.53,    2.53,
  2.94,    2.94,    2.94,    2.94,
  3.13,    3.13,    3.13,    3.13,
  3.11,    3.11,    3.11,    3.11,
  3.48,    3.48,    3.48,    3.48,
  3.64,    3.64,    3.64,    3.64,
  3.92,    3.92,    3.92,    3.92,
  4.49,    4.49,    4.49,    4.49,
  3.92,    3.92,    3.92,    3.92,
  4.53,    4.53,    4.53,    4.53,
  4.95,    4.95,    4.95,    4.95,
  4.09,    4.09,    4.09,    4.09,
  3.79,    3.79,    3.79,    3.79,
  4.09,    4.09,    4.09,    4.09,
  4.26,    4.26,    4.26,    4.26,
  3.93,    3.93,    3.93,    3.93,
  4.06,    4.06,    4.06,    4.06,
  3.05,    3.05,    3.05,    3.05,
  3.63,    3.63,    3.63,    3.63,
  3.88,    3.88,    3.88,    3.88,
  3.39,    3.39,    3.39,    3.39,
  2.39,    2.39,    2.39,    2.39,
  2.44,    2.44,    2.44,    2.44,
  2.18,    2.18,    2.18,    2.18,
  2.13,    2.13,    2.13,    2.13,
  2.14,    2.14,    2.14,    2.14,
  2.13,    2.13,    2.13,    2.13,
  2.31,    2.31,    2.31,    2.31,
  2.26,    2.26,    2.26,    2.26,
  2.29,    2.29,    2.29,    2.29,
  2.19,    2.19,    2.19,    2.19,
  2.19,    2.19,    2.19,    2.19,
  2.39,    2.39,    2.39,    2.39,
  2.31,    2.31,    2.31,    2.31,
  2.22,    2.22,    2.22,    2.22,
  1.76,    1.76,    1.76,    1.76,
  2.46,    2.46,    2.46,    2.46,
  2.47,    2.47,    2.47,    2.47,
  2.28,    2.28,    2.28,    2.28,
  2.22,    2.22,    2.22,    2.22,
  2.11,    2.11,    2.11,    2.11,
  2.19,    2.19,    2.19,    2.19,
  2.04,    2.04,    2.04,    2.04,
  1.9,     1.9,     1.9,     1.9,
  2.25,    2.25,    2.25,    2.25,
  2.12,    2.12,    2.12,    2.12,
  2.28,    2.28,    2.28,    2.28,
  2.38,    2.38,    2.38,    2.38,
  2.24,    2.24,    2.24,    2.24,
  2.18,    2.18,    2.18,    2.18,
  1.76,    1.76,    1.76,    1.76,
  1.85,    1.85,    1.85,    1.85,
  1.84,    1.84,    1.84,    1.84,
  2.48,    2.48,    2.48,    2.48,
  3.38,    3.38,    3.38,    3.38,
  3.45,    3.45,    3.45,    3.45,
  3.65,    3.65,    3.65,    3.65,
  3.84,    3.84,    3.84,    3.84,
  3.73,    3.73,    3.73,    3.73,
  3.64,    3.64,    3.64,    3.64,
  3.78,    3.78,    3.78,    3.78,
  3.52,    3.52,    3.52,    3.52,
  3.81,    3.81,    3.81,    3.81,
  3.34,    3.34,    3.34,    3.34,
  3.17,    3.17,    3.17,    3.17,
  3.53,    3.53,    3.53,    3.53,
  3.12,    3.12,    3.12,    3.12,
  2.61,    2.61,    2.61,    2.61,
  2.07,    2.07,    2.07,    2.07,
  1.72,    1.72,    1.72,    1.72,
  2.25,    2.25,    2.25,    2.25,
  2.24,    2.24,    2.24,    2.24,
  2.21,    2.21,    2.21,    2.21,
  2.24,    2.24,    2.24,    2.24,
  2.46,    2.46,    2.46,    2.46,
  2.51,    2.51,    2.51,    2.51,
  2.27,    2.27,    2.27,    2.27,
  2.47,    2.47,    2.47,    2.47,
  2.55,    2.55,    2.55,    2.55,
  2.62,    2.62,    2.62,    2.62,
  2.91,    2.91,    2.91,    2.91,
  3.06,    3.06,    3.06,    3.06,
  2.81,    2.81,    2.81,    2.81,
  2.53,    2.53,    2.53,    2.53,
  2.36,    2.36,    2.36,    2.36,
  2.47,    2.47,    2.47,    2.47,
  2.19,    2.19,    2.19,    2.19,
  2.5,     2.5,     2.5,     2.5,
  2.72,    2.72,    2.72,    2.72,
  2.27,    2.27,    2.27,    2.27,
  2.5,     2.5,     2.5,     2.5,
  2.32,    2.32,    2.32,    2.32,
  2.43,    2.43,    2.43,    2.43,
  2.22,    2.22,    2.22,    2.22,
  2.16,    2.16,    2.16,    2.16,
  2.23,    2.23,    2.23,    2.23,
  2.16,    2.16,    2.16,    2.16,
  2.13,    2.13,    2.13,    2.13,
  2.26,    2.26,    2.26,    2.26,
  2.02,    2.02,    2.02,    2.02,
  2.61,    2.61,    2.61,    2.61,
  2.36,    2.36,    2.36,    2.36,
  2.81,    2.81,    2.81,    2.81,
  2.12,    2.12,    2.12,    2.12,
  2.34,    2.34,    2.34,    2.34,
  2.31,    2.31,    2.31,    2.31,
  1.83,    1.83,    1.83,    1.83,
  1.41,    1.41,    1.41,    1.41,
  1.21,    1.21,    1.21,    1.21,
  1.37,    1.37,    1.37,    1.37,
  0.8,     0.8,     0.8,     0.8,
  1.37,    1.37,    1.37,    1.37,
  1.01,    1.01,    1.01,    1.01,
  0.83,    0.83,    0.83,    0.83,
  0.69,    0.69,    0.69,    0.69,
  1.57,    1.57,    1.57,    1.57,
  0.89,    0.89,    0.89,    0.89,
  0.83,    0.83,    0.83,    0.83,
  0.79,    0.79,    0.79,    0.79,
  0.88,    0.88,    0.88,    0.88,
  1.21,    1.21,    1.21,    1.21,
  1.27,    1.27,    1.27,    1.27,
  1.3,     1.3,     1.3,     1.3,
  1.24,    1.24,    1.24,    1.24,
  1.28,    1.28,    1.28,    1.28,
  1.7,     1.7,     1.7,     1.7,
  1.67,    1.67,    1.67,    1.67,
  1.26,    1.26,    1.26,    1.26,
  1.51,    1.51,    1.51,    1.51,
  1.75,    1.75,    1.75,    1.75,
  1.57,    1.57,    1.57,    1.57,
  1.83,    1.83,    1.83,    1.83,
  1.49,    1.49,    1.49,    1.49,
  1.9,     1.9,     1.9,     1.9,
  2.06,    2.06,    2.06,    2.06,
  2.11,    2.11,    2.11,    2.11,
  2.19,    2.19,    2.19,    2.19,
  2.23,    2.23,    2.23,    2.23,
  2.42,    2.42,    2.42,    2.42,
  2.07,    2.07,    2.07,    2.07,
  1.94,    1.94,    1.94,    1.94,
  2.04,    2.04,    2.04,    2.04,
  2.42,    2.42,    2.42,    2.42,
  2.5,     2.5,     2.5,     2.5,
  2.48,    2.48,    2.48,    2.48,
  2.3,     2.3,     2.3,     2.3,
  2.4,     2.4,     2.4,     2.4,
  2.62,    2.62,    2.62,    2.62,
  2.38,    2.38,    2.38,    2.38,
  2.44,    2.44,    2.44,    2.44,
  2.19,    2.19,    2.19,    2.19,
  2.21,    2.21,    2.21,    2.21,
  2.71,    2.71,    2.71,    2.71,
  2.22,    2.22,    2.22,    2.22,
  2.22,    2.22,    2.22,    2.22,
  1.96,    1.96,    1.96,    1.96,
  2.08,    2.08,    2.08,    2.08,
  2.12,    2.12,    2.12,    2.12,
  1.93,    1.93,    1.93,    1.93,
  1.85,    1.85,    1.85,    1.85,
  0.99,    0.99,    0.99,    0.99,
  1.78,    1.78,    1.78,    1.78,
  2.4,     2.4,     2.4,     2.4,
  2.68,    2.68,    2.68,    2.68,
  2.86,    2.86,    2.86,    2.86,
  2,       2,       2,       2,
  1.79,    1.79,    1.79,    1.79,
  1.97,    1.97,    1.97,    1.97,
  2.04,    2.04,    2.04,    2.04,
  2.07,    2.07,    2.07,    2.07,
  2.17,    2.17,    2.17,    2.17,
  1.99,    1.99,    1.99,    1.99,
  1.93,    1.93,    1.93,    1.93,
  2.08,    2.08,    2.08,    2.08,
  2.26,    2.26,    2.26,    2.26,
  2.45,    2.45,    2.45,    2.45,
  2.43,    2.43,    2.43,    2.43,
  2.36,    2.36,    2.36,    2.36,
  2.64,    2.64,    2.64,    2.64,
  2.82,    2.82,    2.82,    2.82,
  2.41,    2.41,    2.41,    2.41,
  3.2,     3.2,     3.2,     3.2,
  2.19,    2.19,    2.19,    2.19,
  2.82,    2.82,    2.82,    2.82,
  2.62,    2.62,    2.62,    2.62,
  1.57,    1.57,    1.57,    1.57,
  1.66,    1.66,    1.66,    1.66,
  2,       2,       2,       2,
  1.98,    1.98,    1.98,    1.98,
  1.93,    1.93,    1.93,    1.93,
  2.05,    2.05,    2.05,    2.05,
  2.23,    2.23,    2.23,    2.23,
  2.34,    2.34,    2.34,    2.34,
  2.57,    2.57,    2.57,    2.57,
  2.36,    2.36,    2.36,    2.36,
  2.62,    2.62,    2.62,    2.62,
  2.82,    2.82,    2.82,    2.82,
  3.53,    3.53,    3.53,    3.53,
  3.49,    3.49,    3.49,    3.49,
  3.85,    3.85,    3.85,    3.85,
  3.79,    3.79,    3.79,    3.79,
  3.1,     3.1,     3.1,     3.1,
  3.82,    3.82,    3.82,    3.82,
  4.1,     4.1,     4.1,     4.1,
  3.43,    3.43,    3.43,    3.43,
  3.05,    3.05,    3.05,    3.05,
  2.93,    2.93,    2.93,    2.93,
  2.61,    2.61,    2.61,    2.61,
  2.5,     2.5,     2.5,     2.5,
  2.87,    2.87,    2.87,    2.87,
  3.72,    3.72,    3.72,    3.72,
  3.13,    3.13,    3.13,    3.13,
  3.29,    3.29,    3.29,    3.29,
  2.71,    2.71,    2.71,    2.71,
  2.21,    2.21,    2.21,    2.21,
  2.28,    2.28,    2.28,    2.28,
  2.27,    2.27,    2.27,    2.27,
  2.71,    2.71,    2.71,    2.71,
  3.02,    3.02,    3.02,    3.02,
  2.65,    2.65,    2.65,    2.65,
  1.93,    1.93,    1.93,    1.93,
  2.38,    2.38,    2.38,    2.38,
  2.31,    2.31,    2.31,    2.31,
  2.61,    2.61,    2.61,    2.61,
  2.6,     2.6,     2.6,     2.6,
  2.9,     2.9,     2.9,     2.9,
  2.42,    2.42,    2.42,    2.42,
  2.36,    2.36,    2.36,    2.36,
  2.46,    2.46,    2.46,    2.46,
  2.68,    2.68,    2.68,    2.68,
  2.58,    2.58,    2.58,    2.58,
  2.45,    2.45,    2.45,    2.45,
  2.28,    2.28,    2.28,    2.28,
  1.99,    1.99,    1.99,    1.99,
  1.99,    1.99,    1.99,    1.99,
  1.57,    1.57,    1.57,    1.57,
  1.42,    1.42,    1.42,    1.42,
  0.11,    0.11,    0.11,    0.11,
  1.42,    1.42,    1.42,    1.42,
  1.68,    1.68,    1.68,    1.68,
  1.78,    1.78,    1.78,    1.78,
  1.36,    1.36,    1.36,    1.36,
  1.06,    1.06,    1.06,    1.06,
  1.51,    1.51,    1.51,    1.51,
  1.77,    1.77,    1.77,    1.77,
  1.75,    1.75,    1.75,    1.75,
  1.99,    1.99,    1.99,    1.99,
  2.03,    2.03,    2.03,    2.03,
  2.35,    2.35,    2.35,    2.35,
  2.63,    2.63,    2.63,    2.63,
  3.04,    3.04,    3.04,    3.04,
  3.04,    3.04,    3.04,    3.04,
  2.16,    2.16,    2.16,    2.16,
  2.11,    2.11,    2.11,    2.11,
  2.87,    2.87,    2.87,    2.87,
  2.66,    2.66,    2.66,    2.66,
  2.89,    2.89,    2.89,    2.89,
  2.77,    2.77,    2.77,    2.77,
  3.03,    3.03,    3.03,    3.03,
  2.97,    2.97,    2.97,    2.97,
  2.65,    2.65,    2.65,    2.65,
  2.3,     2.3,     2.3,     2.3,
  2.56,    2.56,    2.56,    2.56,
  2.37,    2.37,    2.37,    2.37,
  2.59,    2.59,    2.59,    2.59,
  2.6,     2.6,     2.6,     2.6,
  2.22,    2.22,    2.22,    2.22,
  2.79,    2.79,    2.79,    2.79,
  2.63,    2.63,    2.63,    2.63,
  2.56,    2.56,    2.56,    2.56,
  2.88,    2.88,    2.88,    2.88,
  2.51,    2.51,    2.51,    2.51,
  2.7,     2.7,     2.7,     2.7,
  2.86,    2.86,    2.86,    2.86,
  3.12,    3.12,    3.12,    3.12,
  3.08,    3.08,    3.08,    3.08,
  2.98,    2.98,    2.98,    2.98,
  2.74,    2.74,    2.74,    2.74,
  2.88,    2.88,    2.88,    2.88,
  2.71,    2.71,    2.71,    2.71,
  2.6,     2.6,     2.6,     2.6,
  2.56,    2.56,    2.56,    2.56,
  2.88,    2.88,    2.88,    2.88,
  2.8,     2.8,     2.8,     2.8,
  2.53,    2.53,    2.53,    2.53,
  2.55,    2.55,    2.55,    2.55,
  2.32,    2.32,    2.32,    2.32,
  2.66,    2.66,    2.66,    2.66,
  2.57,    2.57,    2.57,    2.57,
  2.44,    2.44,    2.44,    2.44,
  2.85,    2.85,    2.85,    2.85,
  3.38,    3.38,    3.38,    3.38,
  3.19,    3.19,    3.19,    3.19,
  3.22,    3.22,    3.22,    3.22,
  2.88,    2.88,    2.88,    2.88,
  3.16,    3.16,    3.16,    3.16,
  3.3,     3.3,     3.3,     3.3,
  3.02,    3.02,    3.02,    3.02,
  3.33,    3.33,    3.33,    3.33,
  3.71,    3.71,    3.71,    3.71,
  2.98,    2.98,    2.98,    2.98,
  2.79,    2.79,    2.79,    2.79,
  3.15,    3.15,    3.15,    3.15,
  3.14,    3.14,    3.14,    3.14,
  2.95,    2.95,    2.95,    2.95,
  3.04,    3.04,    3.04,    3.04,
  2.67,    2.67,    2.67,    2.67,
  2.89,    2.89,    2.89,    2.89,
  2.83,    2.83,    2.83,    2.83,
  2.19,    2.19,    2.19,    2.19,
  1.89,    1.89,    1.89,    1.89,
  1.84,    1.84,    1.84,    1.84,
  2.26,    2.26,    2.26,    2.26,
  2.56,    2.56,    2.56,    2.56,
  2.49,    2.49,    2.49,    2.49,
  2.71,    2.71,    2.71,    2.71,
  2.84,    2.84,    2.84,    2.84,
  2.82,    2.82,    2.82,    2.82,
  3.17,    3.17,    3.17,    3.17,
  3.23,    3.23,    3.23,    3.23,
  3.31,    3.31,    3.31,    3.31,
  3.13,    3.13,    3.13,    3.13,
  2.97,    2.97,    2.97,    2.97,
  2.77,    2.77,    2.77,    2.77,
  3.12,    3.12,    3.12,    3.12,
  3.19,    3.19,    3.19,    3.19,
  3.13,    3.13,    3.13,    3.13,
  3.15,    3.15,    3.15,    3.15,
  3.26,    3.26,    3.26,    3.26,
  2.97,    2.97,    2.97,    2.97,
  2.92,    2.92,    2.92,    2.92,
  2.94,    2.94,    2.94,    2.94,
  2.65,    2.65,    2.65,    2.65,
  2.66,    2.66,    2.66,    2.66,
  2.63,    2.63,    2.63,    2.63,
  2.41,    2.41,    2.41,    2.41,
  2.38,    2.38,    2.38,    2.38,
  2.97,    2.97,    2.97,    2.97,
  3.5,     3.5,     3.5,     3.5,
  3.01,    3.01,    3.01,    3.01,
  2.86,    2.86,    2.86,    2.86,
  2.75,    2.75,    2.75,    2.75,
  2.51,    2.51,    2.51,    2.51,
  2.74,    2.74,    2.74,    2.74,
  2.77,    2.77,    2.77,    2.77,
  3.1,     3.1,     3.1,     3.1,
  2.88,    2.88,    2.88,    2.88,
  2.62,    2.62,    2.62,    2.62,
  2.47,    2.47,    2.47,    2.47,
  2.48,    2.48,    2.48,    2.48,
  2.09,    2.09,    2.09,    2.09,
  2.29,    2.29,    2.29,    2.29,
  2.96,    2.96,    2.96,    2.96,
  2.55,    2.55,    2.55,    2.55,
  2.55,    2.55,    2.55,    2.55,
  2.83,    2.83,    2.83,    2.83,
  2.77,    2.77,    2.77,    2.77,
  2.32,    2.32,    2.32,    2.32,
  2.39,    2.39,    2.39,    2.39,
  2.28,    2.28,    2.28,    2.28,
  2.13,    2.13,    2.13,    2.13,
  2.11,    2.11,    2.11,    2.11,
  2.57,    2.57,    2.57,    2.57,
  2.55,    2.55,    2.55,    2.55,
  2.51,    2.51,    2.51,    2.51,
  2.57,    2.57,    2.57,    2.57,
  3,       3,       3,       3,
  2.7,     2.7,     2.7,     2.7,
  2.37,    2.37,    2.37,    2.37,
  2.3,     2.3,     2.3,     2.3,
  2.53,    2.53,    2.53,    2.53,
  3.1,     3.1,     3.1,     3.1,
  3.12,    3.12,    3.12,    3.12,
  2.88,    2.88,    2.88,    2.88,
  2.95,    2.95,    2.95,    2.95,
  3.02,    3.02,    3.02,    3.02,
  2.79,    2.79,    2.79,    2.79,
  2.53,    2.53,    2.53,    2.53,
  2.04,    2.04,    2.04,    2.04,
  2.01,    2.01,    2.01,    2.01,
  1.95,    1.95,    1.95,    1.95,
  2.08,    2.08,    2.08,    2.08,
  1.99,    1.99,    1.99,    1.99,
  1.73,    1.73,    1.73,    1.73,
  1.81,    1.81,    1.81,    1.81,
  1.15,    1.15,    1.15,    1.15,
  0.77,    0.77,    0.77,    0.77,
  1.16,    1.16,    1.16,    1.16,
  1.56,    1.56,    1.56,    1.56,
  2.24,    2.24,    2.24,    2.24,
  2.98,    2.98,    2.98,    2.98,
  3.27,    3.27,    3.27,    3.27,
  3.36,    3.36,    3.36,    3.36,
  3.46,    3.46,    3.46,    3.46,
  3.01,    3.01,    3.01,    3.01,
  3.03,    3.03,    3.03,    3.03,
  2.49,    2.49,    2.49,    2.49,
  2.95,    2.95,    2.95,    2.95,
  2.88,    2.88,    2.88,    2.88,
  3.17,    3.17,    3.17,    3.17,
  2.94,    2.94,    2.94,    2.94,
  2.8,     2.8,     2.8,     2.8,
  2.97,    2.97,    2.97,    2.97,
  2.16,    2.16,    2.16,    2.16,
  1.98,    1.98,    1.98,    1.98,
  1.7,     1.7,     1.7,     1.7,
  1.55,    1.55,    1.55,    1.55,
  1.6,     1.6,     1.6,     1.6,
  1.46,    1.46,    1.46,    1.46,
  1.43,    1.43,    1.43,    1.43,
  1.46,    1.46,    1.46,    1.46,
  1.26,    1.26,    1.26,    1.26,
  1.06,    1.06,    1.06,    1.06,
  1.24,    1.24,    1.24,    1.24,
  1.34,    1.34,    1.34,    1.34,
  1.68,    1.68,    1.68,    1.68,
  1.75,    1.75,    1.75,    1.75,
  2.06,    2.06,    2.06,    2.06,
  1.97,    1.97,    1.97,    1.97,
  1.6,     1.6,     1.6,     1.6,
  1.37,    1.37,    1.37,    1.37,
  1.61,    1.61,    1.61,    1.61,
  2.16,    2.16,    2.16,    2.16,
  1.86,    1.86,    1.86,    1.86,
  1.89,    1.89,    1.89,    1.89,
  1.09,    1.09,    1.09,    1.09,
  0.84,    0.84,    0.84,    0.84,
  1.16,    1.16,    1.16,    1.16,
  1.13,    1.13,    1.13,    1.13,
  0.82,    0.82,    0.82,    0.82,
  0.24,    0.24,    0.24,    0.24,
  0.18,    0.18,    0.18,    0.18,
  0.65,    0.65,    0.65,    0.65,
  1.01,    1.01,    1.01,    1.01,
  1.05,    1.05,    1.05,    1.05,
  1.2,     1.2,     1.2,     1.2,
  1.05,    1.05,    1.05,    1.05,
  1.32,    1.32,    1.32,    1.32,
  1.53,    1.53,    1.53,    1.53,
  1.72,    1.72,    1.72,    1.72,
  1.33,    1.33,    1.33,    1.33,
  1.56,    1.56,    1.56,    1.56,
  1.39,    1.39,    1.39,    1.39,
  2.2,     2.2,     2.2,     2.2,
  1.89,    1.89,    1.89,    1.89,
  1.77,    1.77,    1.77,    1.77,
  1.82,    1.82,    1.82,    1.82,
  2.07,    2.07,    2.07,    2.07,
  1.66,    1.66,    1.66,    1.66,
  1.69,    1.69,    1.69,    1.69,
  1.41,    1.41,    1.41,    1.41,
  1.84,    1.84,    1.84,    1.84,
  1.49,    1.49,    1.49,    1.49,
  1.17,    1.17,    1.17,    1.17,
  1.35,    1.35,    1.35,    1.35,
  1.67,    1.67,    1.67,    1.67,
  1.7,     1.7,     1.7,     1.7,
  1.66,    1.66,    1.66,    1.66,
  1.63,    1.63,    1.63,    1.63,
  1.78,    1.78,    1.78,    1.78,
  1.72,    1.72,    1.72,    1.72,
  2.05,    2.05,    2.05,    2.05,
  2.34,    2.34,    2.34,    2.34,
  1.97,    1.97,    1.97,    1.97,
  2.3,     2.3,     2.3,     2.3,
  2.06,    2.06,    2.06,    2.06,
  2.27,    2.27,    2.27,    2.27,
  2.71,    2.71,    2.71,    2.71,
  2.87,    2.87,    2.87,    2.87,
  2.95,    2.95,    2.95,    2.95,
  2.86,    2.86,    2.86,    2.86,
  2.7,     2.7,     2.7,     2.7,
  2.6,     2.6,     2.6,     2.6,
  2.82,    2.82,    2.82,    2.82,
  2.92,    2.92,    2.92,    2.92,
  2.71,    2.71,    2.71,    2.71,
  2.62,    2.62,    2.62,    2.62,
  2.96,    2.96,    2.96,    2.96,
  3.18,    3.18,    3.18,    3.18,
  2.93,    2.93,    2.93,    2.93,
  2.45,    2.45,    2.45,    2.45,
  2.24,    2.24,    2.24,    2.24,
  1.64,    1.64,    1.64,    1.64,
  1.78,    1.78,    1.78,    1.78,
  1.78,    1.78,    1.78,    1.78,
  1.29,    1.29,    1.29,    1.29,
  1.71,    1.71,    1.71,    1.71,
  2.06,    2.06,    2.06,    2.06,
  1.81,    1.81,    1.81,    1.81,
  2.25,    2.25,    2.25,    2.25,
  2.3,     2.3,     2.3,     2.3,
  2.04,    2.04,    2.04,    2.04,
  2.4,     2.4,     2.4,     2.4,
  2.76,    2.76,    2.76,    2.76,
  2.69,    2.69,    2.69,    2.69,
  3.05,    3.05,    3.05,    3.05,
  2.73,    2.73,    2.73,    2.73,
  3.48,    3.48,    3.48,    3.48,
  2.37,    2.37,    2.37,    2.37,
  2.71,    2.71,    2.71,    2.71,
  2.4,     2.4,     2.4,     2.4,
  2.09,    2.09,    2.09,    2.09,
  2.32,    2.32,    2.32,    2.32,
  2.42,    2.42,    2.42,    2.42,
  2.35,    2.35,    2.35,    2.35,
  2.98,    2.98,    2.98,    2.98,
  1.91,    1.91,    1.91,    1.91,
  2.34,    2.34,    2.34,    2.34,
  2.49,    2.49,    2.49,    2.49,
  2.45,    2.45,    2.45,    2.45,
  2.87,    2.87,    2.87,    2.87,
  2.88,    2.88,    2.88,    2.88,
  2.43,    2.43,    2.43,    2.43,
  2.65,    2.65,    2.65,    2.65,
  2.66,    2.66,    2.66,    2.66,
  2.51,    2.51,    2.51,    2.51,
  2.6,     2.6,     2.6,     2.6,
  2.66,    2.66,    2.66,    2.66,
  2.3,     2.3,     2.3,     2.3,
  2.24,    2.24,    2.24,    2.24,
  2.48,    2.48,    2.48,    2.48,
  2.5,     2.5,     2.5,     2.5,
  2.52,    2.52,    2.52,    2.52,
  2.6,     2.6,     2.6,     2.6,
  2.34,    2.34,    2.34,    2.34,
  1.95,    1.95,    1.95,    1.95,
  2.52,    2.52,    2.52,    2.52,
  2.56,    2.56,    2.56,    2.56,
  2.56,    2.56,    2.56,    2.56,
  2.42,    2.42,    2.42,    2.42,
  2.42,    2.42,    2.42,    2.42,
  2.81,    2.81,    2.81,    2.81,
  2.59,    2.59,    2.59,    2.59,
  3.4,     3.4,     3.4,     3.4,
  2.8,     2.8,     2.8,     2.8,
  2.66,    2.66,    2.66,    2.66,
  2.87,    2.87,    2.87,    2.87,
  1.91,    1.91,    1.91,    1.91,
  1.88,    1.88,    1.88,    1.88,
  2.51,    2.51,    2.51,    2.51,
  1.97,    1.97,    1.97,    1.97,
  1.95,    1.95,    1.95,    1.95,
  1.94,    1.94,    1.94,    1.94,
  2.01,    2.01,    2.01,    2.01,
  1.82,    1.82,    1.82,    1.82,
  1.87,    1.87,    1.87,    1.87,
  2.51,    2.51,    2.51,    2.51,
  2.63,    2.63,    2.63,    2.63,
  2.51,    2.51,    2.51,    2.51,
  2.04,    2.04,    2.04,    2.04,
  2.07,    2.07,    2.07,    2.07,
  2.19,    2.19,    2.19,    2.19,
  2.29,    2.29,    2.29,    2.29,
  2.62,    2.62,    2.62,    2.62,
  2.31,    2.31,    2.31,    2.31,
  2.47,    2.47,    2.47,    2.47,
  2.5,     2.5,     2.5,     2.5,
  2.38,    2.38,    2.38,    2.38,
  2.57,    2.57,    2.57,    2.57,
  2.68,    2.68,    2.68,    2.68,
  2.84,    2.84,    2.84,    2.84,
  2.77,    2.77,    2.77,    2.77,
  2.38,    2.38,    2.38,    2.38,
  2.42,    2.42,    2.42,    2.42,
  2.69,    2.69,    2.69,    2.69,
  2.83,    2.83,    2.83,    2.83,
  2.36,    2.36,    2.36,    2.36,
  1.81,    1.81,    1.81,    1.81,
  1.46,    1.46,    1.46,    1.46,
  1.7,     1.7,     1.7,     1.7,
  1.47,    1.47,    1.47,    1.47,
  1.48,    1.48,    1.48,    1.48,
  1.55,    1.55,    1.55,    1.55,
  1.55,    1.55,    1.55,    1.55,
  1.3,     1.3,     1.3,     1.3,
  1.14,    1.14,    1.14,    1.14,
  1.65,    1.65,    1.65,    1.65,
  2,       2,       2,       2,
  2.58,    2.58,    2.58,    2.58,
  2.35,    2.35,    2.35,    2.35,
  2.45,    2.45,    2.45,    2.45,
  2.31,    2.31,    2.31,    2.31,
  2.25,    2.25,    2.25,    2.25,
  1.85,    1.85,    1.85,    1.85,
  2.36,    2.36,    2.36,    2.36,
  2.31,    2.31,    2.31,    2.31,
  2.04,    2.04,    2.04,    2.04,
  1.38,    1.38,    1.38,    1.38,
  1.19,    1.19,    1.19,    1.19,
  1.3,     1.3,     1.3,     1.3,
  1.32,    1.32,    1.32,    1.32,
  1.71,    1.71,    1.71,    1.71,
  1.54,    1.54,    1.54,    1.54,
  1.71,    1.71,    1.71,    1.71,
  1.88,    1.88,    1.88,    1.88,
  1.25,    1.25,    1.25,    1.25,
  1.26,    1.26,    1.26,    1.26,
  0.96,    0.96,    0.96,    0.96,
  1.07,    1.07,    1.07,    1.07,
  1.87,    1.87,    1.87,    1.87,
  1.91,    1.91,    1.91,    1.91,
  2.15,    2.15,    2.15,    2.15,
  3.01,    3.01,    3.01,    3.01,
  2.64,    2.64,    2.64,    2.64,
  2.08,    2.08,    2.08,    2.08,
  2.23,    2.23,    2.23,    2.23,
  2.5,     2.5,     2.5,     2.5,
  2.21,    2.21,    2.21,    2.21,
  1.48,    1.48,    1.48,    1.48,
  1.71,    1.71,    1.71,    1.71,
  1.98,    1.98,    1.98,    1.98,
  1.79,    1.79,    1.79,    1.79,
  1.7,     1.7,     1.7,     1.7,
  1.71,    1.71,    1.71,    1.71,
  2.04,    2.04,    2.04,    2.04,
  1.63,    1.63,    1.63,    1.63,
  1.9,     1.9,     1.9,     1.9,
  1.73,    1.73,    1.73,    1.73,
  1.45,    1.45,    1.45,    1.45,
  1.54,    1.54,    1.54,    1.54,
  1.42,    1.42,    1.42,    1.42,
  0.97,    0.97,    0.97,    0.97,
  0.87,    0.87,    0.87,    0.87,
  0.95,    0.95,    0.95,    0.95,
  0.72,    0.72,    0.72,    0.72,
  0.75,    0.75,    0.75,    0.75,
  0.62,    0.62,    0.62,    0.62,
  0.51,    0.51,    0.51,    0.51,
  0.63,    0.63,    0.63,    0.63,
  0.46,    0.46,    0.46,    0.46,
  0.42,    0.42,    0.42,    0.42,
  0.62,    0.62,    0.62,    0.62,
  0.91,    0.91,    0.91,    0.91,
  0.67,    0.67,    0.67,    0.67,
  0.48,    0.48,    0.48,    0.48,
  0.63,    0.63,    0.63,    0.63,
  1.25,    1.25,    1.25,    1.25,
  1.56,    1.56,    1.56,    1.56,
  1.36,    1.36,    1.36,    1.36,
  1.22,    1.22,    1.22,    1.22,
  1.28,    1.28,    1.28,    1.28,
  1.36,    1.36,    1.36,    1.36,
  2.03,    2.03,    2.03,    2.03,
  1.86,    1.86,    1.86,    1.86,
  1.4,     1.4,     1.4,     1.4,
  1.37,    1.37,    1.37,    1.37,
  1.64,    1.64,    1.64,    1.64,
  1.42,    1.42,    1.42,    1.42,
  1.24,    1.24,    1.24,    1.24,
  1.47,    1.47,    1.47,    1.47,
  1.48,    1.48,    1.48,    1.48,
  1.21,    1.21,    1.21,    1.21,
  1.02,    1.02,    1.02,    1.02,
  0.92,    0.92,    0.92,    0.92,
  1.32,    1.32,    1.32,    1.32,
  1.85,    1.85,    1.85,    1.85,
  1.18,    1.18,    1.18,    1.18,
  1.46,    1.46,    1.46,    1.46,
  1.49,    1.49,    1.49,    1.49,
  0.96,    0.96,    0.96,    0.96,
  1.25,    1.25,    1.25,    1.25,
  1.61,    1.61,    1.61,    1.61,
  1.82,    1.82,    1.82,    1.82,
  1.48,    1.48,    1.48,    1.48,
  0.75,    0.75,    0.75,    0.75,
  1.64,    1.64,    1.64,    1.64,
  1.21,    1.21,    1.21,    1.21,
  1.3,     1.3,     1.3,     1.3,
  1.37,    1.37,    1.37,    1.37,
  0.77,    0.77,    0.77,    0.77,
  1.28,    1.28,    1.28,    1.28,
  1.1,     1.1,     1.1,     1.1,
  0.24,    0.24,    0.24,    0.24,
  0.82,    0.82,    0.82,    0.82,
  0.4,     0.4,     0.4,     0.4,
  1.35,    1.35,    1.35,    1.35,
  0.64,    0.64,    0.64,    0.64,
  0.64,    0.64,    0.64,    0.64,
  0.79,    0.79,    0.79,    0.79,
  0.7,     0.7,     0.7,     0.7,
  0.83,    0.83,    0.83,    0.83,
  1.07,    1.07,    1.07,    1.07,
  1.24,    1.24,    1.24,    1.24,
  1.55,    1.55,    1.55,    1.55,
  1.19,    1.19,    1.19,    1.19,
  1.65,    1.65,    1.65,    1.65,
  1.91,    1.91,    1.91,    1.91,
  1.69,    1.69,    1.69,    1.69,
  1.86,    1.86,    1.86,    1.86,
  1.74,    1.74,    1.74,    1.74,
  1.19,    1.19,    1.19,    1.19,
  1,       1,       1,       1,
  0.66,    0.66,    0.66,    0.66,
  1.23,    1.23,    1.23,    1.23,
  0.95,    0.95,    0.95,    0.95,
  1.02,    1.02,    1.02,    1.02,
  1.73,    1.73,    1.73,    1.73,
  1.83,    1.83,    1.83,    1.83,
  1.43,    1.43,    1.43,    1.43,
  1.02,    1.02,    1.02,    1.02,
  0.78,    0.78,    0.78,    0.78,
  1,       1,       1,       1,
  1.06,    1.06,    1.06,    1.06,
  1.16,    1.16,    1.16,    1.16,
  1.51,    1.51,    1.51,    1.51,
  0.98,    0.98,    0.98,    0.98,
  0.99,    0.99,    0.99,    0.99,
  1.12,    1.12,    1.12,    1.12,
  0.78,    0.78,    0.78,    0.78,
  1.02,    1.02,    1.02,    1.02,
  1.29,    1.29,    1.29,    1.29,
  1.69,    1.69,    1.69,    1.69,
  1.11,    1.11,    1.11,    1.11,
  1,       1,       1,       1,
  0.91,    0.91,    0.91,    0.91,
  1.21,    1.21,    1.21,    1.21,
  1.05,    1.05,    1.05,    1.05,
  0.81,    0.81,    0.81,    0.81,
  0.37,    0.37,    0.37,    0.37,
  0.36,    0.36,    0.36,    0.36,
  0.49,    0.49,    0.49,    0.49,
  0.52,    0.52,    0.52,    0.52,
  0.94,    0.94,    0.94,    0.94,
  1.16,    1.16,    1.16,    1.16,
  1.17,    1.17,    1.17,    1.17,
  1.21,    1.21,    1.21,    1.21,
  1.13,    1.13,    1.13,    1.13,
  1.06,    1.06,    1.06,    1.06,
  0.87,    0.87,    0.87,    0.87,
  0.81,    0.81,    0.81,    0.81,
  0.95,    0.95,    0.95,    0.95,
  1.56,    1.56,    1.56,    1.56,
  1.12,    1.12,    1.12,    1.12,
  0.91,    0.91,    0.91,    0.91,
  0.88,    0.88,    0.88,    0.88,
  0.23,    0.23,    0.23,    0.23,
  0.75,    0.75,    0.75,    0.75,
  0.91,    0.91,    0.91,    0.91,
  1.07,    1.07,    1.07,    1.07,
  0.28,    0.28,    0.28,    0.28,
  1.02,    1.02,    1.02,    1.02,
  0.78,    0.78,    0.78,    0.78,
  1.3,     1.3,     1.3,     1.3,
  0.29,    0.29,    0.29,    0.29,
  0.37,    0.37,    0.37,    0.37,
  1.06,    1.06,    1.06,    1.06,
  1.08,    1.08,    1.08,    1.08,
  0.37,    0.37,    0.37,    0.37,
  1.4,     1.4,     1.4,     1.4,
  2.36,    2.36,    2.36,    2.36,
  2.84,    2.84,    2.84,    2.84,
  2.81,    2.81,    2.81,    2.81,
  2.72,    2.72,    2.72,    2.72,
  2.59,    2.59,    2.59,    2.59,
  1.74,    1.74,    1.74,    1.74,
  1.74,    1.74,    1.74,    1.74,
  2.17,    2.17,    2.17,    2.17,
  2.17,    2.17,    2.17,    2.17,
  2.03,    2.03,    2.03,    2.03,
  1.56,    1.56,    1.56,    1.56,
  2.18,    2.18,    2.18,    2.18,
  0.88,    0.88,    0.88,    0.88,
  0.95,    0.95,    0.95,    0.95,
  0.43,    0.43,    0.43,    0.43,
  0.98,    0.98,    0.98,    0.98,
  0.5,     0.5,     0.5,     0.5,
  0.26,    0.26,    0.26,    0.26,
  0.39,    0.39,    0.39,    0.39,
  0.9,     0.9,     0.9,     0.9,
  1.8,     1.8,     1.8,     1.8,
  2.21,    2.21,    2.21,    2.21,
  2.66,    2.66,    2.66,    2.66,
  2.48,    2.48,    2.48,    2.48,
  2.4,     2.4,     2.4,     2.4,
  2.54,    2.54,    2.54,    2.54,
  2.97,    2.97,    2.97,    2.97,
  3.28,    3.28,    3.28,    3.28,
  4.06,    4.06,    4.06,    4.06,
  4.06,    4.06,    4.06,    4.06,
  3.7,     3.7,     3.7,     3.7,
  4.29,    4.29,    4.29,    4.29,
  3.9,     3.9,     3.9,     3.9,
  4.2,     4.2,     4.2,     4.2,
  3.95,    3.95,    3.95,    3.95,
  4.44,    4.44,    4.44,    4.44,
  4.2,     4.2,     4.2,     4.2,
  4.48,    4.48,    4.48,    4.48,
  3.36,    3.36,    3.36,    3.36,
  3,       3,       3,       3,
  2.87,    2.87,    2.87,    2.87,
  3.17,    3.17,    3.17,    3.17,
  3.86,    3.86,    3.86,    3.86,
  3.49,    3.49,    3.49,    3.49,
  3.92,    3.92,    3.92,    3.92,
  3.83,    3.83,    3.83,    3.83,
  4.29,    4.29,    4.29,    4.29,
  4,       4,       4,       4,
  3.91,    3.91,    3.91,    3.91,
  4.01,    4.01,    4.01,    4.01,
  3.84,    3.84,    3.84,    3.84,
  2.92,    2.92,    2.92,    2.92,
  3.84,    3.84,    3.84,    3.84,
  3.45,    3.45,    3.45,    3.45,
  4.1,     4.1,     4.1,     4.1,
  3.87,    3.87,    3.87,    3.87,
  3.67,    3.67,    3.67,    3.67,
  3.55,    3.55,    3.55,    3.55,
  4.03,    4.03,    4.03,    4.03,
  3.75,    3.75,    3.75,    3.75,
  3.75,    3.75,    3.75,    3.75,
  3.63,    3.63,    3.63,    3.63,
  3.47,    3.47,    3.47,    3.47,
  3.34,    3.34,    3.34,    3.34,
  2.79,    2.79,    2.79,    2.79,
  3.35,    3.35,    3.35,    3.35,
  3.36,    3.36,    3.36,    3.36,
  3.19,    3.19,    3.19,    3.19,
  3.72,    3.72,    3.72,    3.72,
  3.6,     3.6,     3.6,     3.6,
  3.45,    3.45,    3.45,    3.45,
  4.58,    4.58,    4.58,    4.58,
  3.95,    3.95,    3.95,    3.95,
  5.37,    5.37,    5.37,    5.37,
  4.69,    4.69,    4.69,    4.69,
  4.27,    4.27,    4.27,    4.27,
  4.83,    4.83,    4.83,    4.83,
  4.52,    4.52,    4.52,    4.52,
  5.4,     5.4,     5.4,     5.4,
  4.53,    4.53,    4.53,    4.53,
  5.2,     5.2,     5.2,     5.2,
  5.12,    5.12,    5.12,    5.12,
  5.04,    5.04,    5.04,    5.04,
  4.32,    4.32,    4.32,    4.32,
  4.73,    4.73,    4.73,    4.73,
  4.7,     4.7,     4.7,     4.7,
  4.4,     4.4,     4.4,     4.4,
  4.94,    4.94,    4.94,    4.94,
  4.02,    4.02,    4.02,    4.02,
  4.13,    4.13,    4.13,    4.13,
  3.8,     3.8,     3.8,     3.8,
  3.16,    3.16,    3.16,    3.16,
  2.75,    2.75,    2.75,    2.75,
  2.51,    2.51,    2.51,    2.51,
  2.85,    2.85,    2.85,    2.85,
  2.87,    2.87,    2.87,    2.87,
  2.56,    2.56,    2.56,    2.56,
  2.38,    2.38,    2.38,    2.38,
  2,       2,       2,       2,
  1.81,    1.81,    1.81,    1.81,
  0.71,    0.71,    0.71,    0.71,
  1.39,    1.39,    1.39,    1.39,
  2.07,    2.07,    2.07,    2.07,
  1.84,    1.84,    1.84,    1.84,
  2.17,    2.17,    2.17,    2.17,
  1.93,    1.93,    1.93,    1.93,
  2.08,    2.08,    2.08,    2.08,
  2.12,    2.12,    2.12,    2.12,
  1.99,    1.99,    1.99,    1.99,
  1.74,    1.74,    1.74,    1.74,
  1.32,    1.32,    1.32,    1.32,
  1.88,    1.88,    1.88,    1.88,
  2.07,    2.07,    2.07,    2.07,
  1.85,    1.85,    1.85,    1.85,
  2.03,    2.03,    2.03,    2.03,
  1.97,    1.97,    1.97,    1.97,
  1.89,    1.89,    1.89,    1.89,
  1.61,    1.61,    1.61,    1.61,
  1.62,    1.62,    1.62,    1.62,
  1.62,    1.62,    1.62,    1.62,
  2.03,    2.03,    2.03,    2.03,
  2.24,    2.24,    2.24,    2.24,
  2.43,    2.43,    2.43,    2.43,
  2.24,    2.24,    2.24,    2.24,
  1.75,    1.75,    1.75,    1.75,
  1.8,     1.8,     1.8,     1.8,
  1.89,    1.89,    1.89,    1.89,
  1.87,    1.87,    1.87,    1.87,
  1.77,    1.77,    1.77,    1.77,
  2.13,    2.13,    2.13,    2.13,
  2.3,     2.3,     2.3,     2.3,
  1.67,    1.67,    1.67,    1.67,
  2.65,    2.65,    2.65,    2.65,
  2,       2,       2,       2,
  1.33,    1.33,    1.33,    1.33,
  1.33,    1.33,    1.33,    1.33,
  1.53,    1.53,    1.53,    1.53,
  1.6,     1.6,     1.6,     1.6,
  2.47,    2.47,    2.47,    2.47,
  2.59,    2.59,    2.59,    2.59,
  2.37,    2.37,    2.37,    2.37,
  2.74,    2.74,    2.74,    2.74,
  2.44,    2.44,    2.44,    2.44,
  2.32,    2.32,    2.32,    2.32,
  2.38,    2.38,    2.38,    2.38,
  2.48,    2.48,    2.48,    2.48,
  2.51,    2.51,    2.51,    2.51,
  2.64,    2.64,    2.64,    2.64,
  2.66,    2.66,    2.66,    2.66,
  2.6,     2.6,     2.6,     2.6,
  2.44,    2.44,    2.44,    2.44,
  2.28,    2.28,    2.28,    2.28,
  1.97,    1.97,    1.97,    1.97,
  2.34,    2.34,    2.34,    2.34,
  2.46,    2.46,    2.46,    2.46,
  2.37,    2.37,    2.37,    2.37,
  2.35,    2.35,    2.35,    2.35,
  2.62,    2.62,    2.62,    2.62,
  2.58,    2.58,    2.58,    2.58,
  2.3,     2.3,     2.3,     2.3,
  2.62,    2.62,    2.62,    2.62,
  2.75,    2.75,    2.75,    2.75,
  2.76,    2.76,    2.76,    2.76,
  2.59,    2.59,    2.59,    2.59,
  2.81,    2.81,    2.81,    2.81,
  2.35,    2.35,    2.35,    2.35,
  2.52,    2.52,    2.52,    2.52,
  2.33,    2.33,    2.33,    2.33,
  2.94,    2.94,    2.94,    2.94,
  2.46,    2.46,    2.46,    2.46,
  2.72,    2.72,    2.72,    2.72,
  3.35,    3.35,    3.35,    3.35,
  3.43,    3.43,    3.43,    3.43,
  3.62,    3.62,    3.62,    3.62,
  3.54,    3.54,    3.54,    3.54,
  3.36,    3.36,    3.36,    3.36,
  3.52,    3.52,    3.52,    3.52,
  3.68,    3.68,    3.68,    3.68,
  2.92,    2.92,    2.92,    2.92,
  3.02,    3.02,    3.02,    3.02,
  3.38,    3.38,    3.38,    3.38,
  2.83,    2.83,    2.83,    2.83,
  3.05,    3.05,    3.05,    3.05,
  3.02,    3.02,    3.02,    3.02,
  2.9,     2.9,     2.9,     2.9,
  2.81,    2.81,    2.81,    2.81,
  2.49,    2.49,    2.49,    2.49,
  2.6,     2.6,     2.6,     2.6,
  2.47,    2.47,    2.47,    2.47,
  2.69,    2.69,    2.69,    2.69,
  2.91,    2.91,    2.91,    2.91,
  2.91,    2.91,    2.91,    2.91,
  2.72,    2.72,    2.72,    2.72,
  2.41,    2.41,    2.41,    2.41,
  2.34,    2.34,    2.34,    2.34,
  2.69,    2.69,    2.69,    2.69,
  2.64,    2.64,    2.64,    2.64,
  2.92,    2.92,    2.92,    2.92,
  2.97,    2.97,    2.97,    2.97,
  2.82,    2.82,    2.82,    2.82,
  2.43,    2.43,    2.43,    2.43,
  2.39,    2.39,    2.39,    2.39,
  2.04,    2.04,    2.04,    2.04,
  2.03,    2.03,    2.03,    2.03,
  2.16,    2.16,    2.16,    2.16,
  2.81,    2.81,    2.81,    2.81,
  2.6,     2.6,     2.6,     2.6,
  2.5,     2.5,     2.5,     2.5,
  2.24,    2.24,    2.24,    2.24,
  2.05,    2.05,    2.05,    2.05,
  1.92,    1.92,    1.92,    1.92,
  2.25,    2.25,    2.25,    2.25,
  2.61,    2.61,    2.61,    2.61,
  2.29,    2.29,    2.29,    2.29,
  1.87,    1.87,    1.87,    1.87,
  2.33,    2.33,    2.33,    2.33,
  1.84,    1.84,    1.84,    1.84,
  1.99,    1.99,    1.99,    1.99,
  1.68,    1.68,    1.68,    1.68,
  1.98,    1.98,    1.98,    1.98,
  2.14,    2.14,    2.14,    2.14,
  2.4,     2.4,     2.4,     2.4,
  2.33,    2.33,    2.33,    2.33,
  2.65,    2.65,    2.65,    2.65,
  2.76,    2.76,    2.76,    2.76,
  2.38,    2.38,    2.38,    2.38,
  2.22,    2.22,    2.22,    2.22,
  2.19,    2.19,    2.19,    2.19,
  2.81,    2.81,    2.81,    2.81,
  2.04,    2.04,    2.04,    2.04,
  1.97,    1.97,    1.97,    1.97,
  1.76,    1.76,    1.76,    1.76,
  1.49,    1.49,    1.49,    1.49,
  1.22,    1.22,    1.22,    1.22,
  1.04,    1.04,    1.04,    1.04,
  1.18,    1.18,    1.18,    1.18,
  1.29,    1.29,    1.29,    1.29,
  1.37,    1.37,    1.37,    1.37,
  1.33,    1.33,    1.33,    1.33,
  1.07,    1.07,    1.07,    1.07,
  1.23,    1.23,    1.23,    1.23,
  1.15,    1.15,    1.15,    1.15,
  1.24,    1.24,    1.24,    1.24,
  1.22,    1.22,    1.22,    1.22,
  1.39,    1.39,    1.39,    1.39,
  1.33,    1.33,    1.33,    1.33,
  1.33,    1.33,    1.33,    1.33,
  1.23,    1.23,    1.23,    1.23,
  1.37,    1.37,    1.37,    1.37,
  1.36,    1.36,    1.36,    1.36,
  1.25,    1.25,    1.25,    1.25,
  1.68,    1.68,    1.68,    1.68,
  1.86,    1.86,    1.86,    1.86,
  2.09,    2.09,    2.09,    2.09,
  2.16,    2.16,    2.16,    2.16,
  2.02,    2.02,    2.02,    2.02,
  2.01,    2.01,    2.01,    2.01,
  2.11,    2.11,    2.11,    2.11,
  1.99,    1.99,    1.99,    1.99,
  1.72,    1.72,    1.72,    1.72,
  1.77,    1.77,    1.77,    1.77,
  1.51,    1.51,    1.51,    1.51,
  1.94,    1.94,    1.94,    1.94,
  1.79,    1.79,    1.79,    1.79,
  2.13,    2.13,    2.13,    2.13,
  2.66,    2.66,    2.66,    2.66,
  2.34,    2.34,    2.34,    2.34,
  2.41,    2.41,    2.41,    2.41,
  2.71,    2.71,    2.71,    2.71,
  3.08,    3.08,    3.08,    3.08,
  3.18,    3.18,    3.18,    3.18,
  3.01,    3.01,    3.01,    3.01,
  2.85,    2.85,    2.85,    2.85,
  2.64,    2.64,    2.64,    2.64,
  2.58,    2.58,    2.58,    2.58,
  2.99,    2.99,    2.99,    2.99,
  2.74,    2.74,    2.74,    2.74,
  2.39,    2.39,    2.39,    2.39,
  1.73,    1.73,    1.73,    1.73,
  1.95,    1.95,    1.95,    1.95,
  2.35,    2.35,    2.35,    2.35,
  2.54,    2.54,    2.54,    2.54,
  2.69,    2.69,    2.69,    2.69,
  2.88,    2.88,    2.88,    2.88,
  2.81,    2.81,    2.81,    2.81,
  2.87,    2.87,    2.87,    2.87,
  2.51,    2.51,    2.51,    2.51,
  2.59,    2.59,    2.59,    2.59,
  2.65,    2.65,    2.65,    2.65,
  2.44,    2.44,    2.44,    2.44,
  2.61,    2.61,    2.61,    2.61,
  2.71,    2.71,    2.71,    2.71,
  2.74,    2.74,    2.74,    2.74,
  2.58,    2.58,    2.58,    2.58,
  2.4,     2.4,     2.4,     2.4,
  2.42,    2.42,    2.42,    2.42,
  3.34,    3.34,    3.34,    3.34,
  2.81,    2.81,    2.81,    2.81,
  1.17,    1.17,    1.17,    1.17,
  2.04,    2.04,    2.04,    2.04,
  2.44,    2.44,    2.44,    2.44,
  2.61,    2.61,    2.61,    2.61,
  2.49,    2.49,    2.49,    2.49,
  2.88,    2.88,    2.88,    2.88,
  2.73,    2.73,    2.73,    2.73,
  2.97,    2.97,    2.97,    2.97,
  3.22,    3.22,    3.22,    3.22,
  3.25,    3.25,    3.25,    3.25,
  3.44,    3.44,    3.44,    3.44,
  3.55,    3.55,    3.55,    3.55,
  3.17,    3.17,    3.17,    3.17,
  3.37,    3.37,    3.37,    3.37,
  3.52,    3.52,    3.52,    3.52,
  3.99,    3.99,    3.99,    3.99,
  4.01,    4.01,    4.01,    4.01,
  4.57,    4.57,    4.57,    4.57,
  5.06,    5.06,    5.06,    5.06,
  5.5,     5.5,     5.5,     5.5,
  6.16,    6.16,    6.16,    6.16,
  2.363,   2.363,   2.363,   2.363,
  2.454,   2.454,   2.454,   2.454,
  2.467,   2.467,   2.467,   2.467,
  2.384,   2.384,   2.384,   2.384,
  2.328,   2.328,   2.328,   2.328,
  4.4,     4.4,     4.4,     4.4,
  3.43,    3.43,    3.43,    3.43,
  3.3,     3.3,     3.3,     3.3,
  3.49,    3.49,    3.49,    3.49,
  3.51,    3.51,    3.51,    3.51,
  3.81,    3.81,    3.81,    3.81,
  3.48,    3.48,    3.48,    3.48,
  3.36,    3.36,    3.36,    3.36,
  3.81,    3.81,    3.81,    3.81,
  3.59,    3.59,    3.59,    3.59,
  3.95,    3.95,    3.95,    3.95,
  3.53,    3.53,    3.53,    3.53,
  3.76,    3.76,    3.76,    3.76,
  3.93,    3.93,    3.93,    3.93,
  3.68,    3.68,    3.68,    3.68,
  3.42,    3.42,    3.42,    3.42,
  3.57,    3.57,    3.57,    3.57,
  3.34,    3.34,    3.34,    3.34,
  3.52,    3.52,    3.52,    3.52,
  3.32,    3.32,    3.32,    3.32,
  3.5,     3.5,     3.5,     3.5,
  3.42,    3.42,    3.42,    3.42,
  3.14,    3.14,    3.14,    3.14,
  3.07,    3.07,    3.07,    3.07,
  3.16,    3.16,    3.16,    3.16,
  3.03,    3.03,    3.03,    3.03,
  3.23,    3.23,    3.23,    3.23,
  3.47,    3.47,    3.47,    3.47,
  3.62,    3.62,    3.62,    3.62,
  3.66,    3.66,    3.66,    3.66,
  4.04,    4.04,    4.04,    4.04,
  3.9,     3.9,     3.9,     3.9,
  3.67,    3.67,    3.67,    3.67,
  3.67,    3.67,    3.67,    3.67,
  3.68,    3.68,    3.68,    3.68,
  4.11,    4.11,    4.11,    4.11,
  3.22,    3.22,    3.22,    3.22,
  3.65,    3.65,    3.65,    3.65,
  3.7,     3.7,     3.7,     3.7,
  3.88,    3.88,    3.88,    3.88,
  4.67,    4.67,    4.67,    4.67,
  4.54,    4.54,    4.54,    4.54,
  4.74,    4.74,    4.74,    4.74,
  4.66,    4.66,    4.66,    4.66,
  4.72,    4.72,    4.72,    4.72,
  5.26,    5.26,    5.26,    5.26,
  5.47,    5.47,    5.47,    5.47,
  4.44,    4.44,    4.44,    4.44,
  4.34,    4.34,    4.34,    4.34,
  4.97,    4.97,    4.97,    4.97,
  5.22,    5.22,    5.22,    5.22,
  4.33,    4.33,    4.33,    4.33,
  4.64,    4.64,    4.64,    4.64,
  5.34,    5.34,    5.34,    5.34,
  5.07,    5.07,    5.07,    5.07,
  5.74,    5.74,    5.74,    5.74,
  6.39,    6.39,    6.39,    6.39,
  6.51,    6.51,    6.51,    6.51,
  6.01,    6.01,    6.01,    6.01,
  6.65,    6.65,    6.65,    6.65,
  6.55,    6.55,    6.55,    6.55,
  6.42,    6.42,    6.42,    6.42,
  5.93,    5.93,    5.93,    5.93,
  6.11,    6.11,    6.11,    6.11,
  6.35,    6.35,    6.35,    6.35,
  6.22,    6.22,    6.22,    6.22,
  5.7,     5.7,     5.7,     5.7,
  5.06,    5.06,    5.06,    5.06,
  4.03,    4.03,    4.03,    4.03,
  3.48,    3.48,    3.48,    3.48,
  2.46,    2.46,    2.46,    2.46,
  3.26,    3.26,    3.26,    3.26,
  3.84,    3.84,    3.84,    3.84,
  4.95,    4.95,    4.95,    4.95,
  4.65,    4.65,    4.65,    4.65,
  5.09,    5.09,    5.09,    5.09,
  5.31,    5.31,    5.31,    5.31,
  5.69,    5.69,    5.69,    5.69,
  5.85,    5.85,    5.85,    5.85,
  5.94,    5.94,    5.94,    5.94,
  5.42,    5.42,    5.42,    5.42,
  5.63,    5.63,    5.63,    5.63,
  6.37,    6.37,    6.37,    6.37,
  6.98,    6.98,    6.98,    6.98,
  7.16,    7.16,    7.16,    7.16,
  6.57,    6.57,    6.57,    6.57,
  6.68,    6.68,    6.68,    6.68,
  6.73,    6.73,    6.73,    6.73,
  7.07,    7.07,    7.07,    7.07,
  6.63,    6.63,    6.63,    6.63,
  6.1,     6.1,     6.1,     6.1,
  5.28,    5.28,    5.28,    5.28,
  7.82,    7.82,    7.82,    7.82,
  6.51,    6.51,    6.51,    6.51,
  6.1,     6.1,     6.1,     6.1,
  6.55,    6.55,    6.55,    6.55,
  5.66,    5.66,    5.66,    5.66,
  5.64,    5.64,    5.64,    5.64,
  6.12,    6.12,    6.12,    6.12,
  6.47,    6.47,    6.47,    6.47,
  6.07,    6.07,    6.07,    6.07,
  5.53,    5.53,    5.53,    5.53,
  4.6,     4.6,     4.6,     4.6,
  4.4,     4.4,     4.4,     4.4,
  4.6,     4.6,     4.6,     4.6,
  4.32,    4.32,    4.32,    4.32,
  3.9,     3.9,     3.9,     3.9,
  3.85,    3.85,    3.85,    3.85,
  3.17,    3.17,    3.17,    3.17,
  3.59,    3.59,    3.59,    3.59,
  3.39,    3.39,    3.39,    3.39,
  2.88,    2.88,    2.88,    2.88,
  3.09,    3.09,    3.09,    3.09,
  3.58,    3.58,    3.58,    3.58,
  3.36,    3.36,    3.36,    3.36,
  3.91,    3.91,    3.91,    3.91,
  4.9,     4.9,     4.9,     4.9,
  5.4,     5.4,     5.4,     5.4,
  5.35,    5.35,    5.35,    5.35,
  5.11,    5.11,    5.11,    5.11,
  3.98,    3.98,    3.98,    3.98,
  4.87,    4.87,    4.87,    4.87,
  3.81,    3.81,    3.81,    3.81,
  4.11,    4.11,    4.11,    4.11,
  3.93,    3.93,    3.93,    3.93,
  3.45,    3.45,    3.45,    3.45,
  4.08,    4.08,    4.08,    4.08,
  5.67,    5.67,    5.67,    5.67,
  4.45,    4.45,    4.45,    4.45,
  4.33,    4.33,    4.33,    4.33,
  5.51,    5.51,    5.51,    5.51,
  6.33,    6.33,    6.33,    6.33,
  5.65,    5.65,    5.65,    5.65,
  6.1,     6.1,     6.1,     6.1,
  6.46,    6.46,    6.46,    6.46,
  6.27,    6.27,    6.27,    6.27,
  6.13,    6.13,    6.13,    6.13,
  6.11,    6.11,    6.11,    6.11,
  6.49,    6.49,    6.49,    6.49,
  6.18,    6.18,    6.18,    6.18,
  6.67,    6.67,    6.67,    6.67,
  5.93,    5.93,    5.93,    5.93,
  6.46,    6.46,    6.46,    6.46,
  6.45,    6.45,    6.45,    6.45,
  6.8,     6.8,     6.8,     6.8,
  6.13,    6.13,    6.13,    6.13,
  5.84,    5.84,    5.84,    5.84,
  5.12,    5.12,    5.12,    5.12,
  4.85,    4.85,    4.85,    4.85,
  3.45,    3.45,    3.45,    3.45,
  4.48,    4.48,    4.48,    4.48,
  4.97,    4.97,    4.97,    4.97,
  3.77,    3.77,    3.77,    3.77,
  4.95,    4.95,    4.95,    4.95,
  5.07,    5.07,    5.07,    5.07,
  4.6,     4.6,     4.6,     4.6,
  4.25,    4.25,    4.25,    4.25,
  3.21,    3.21,    3.21,    3.21,
  2.35,    2.35,    2.35,    2.35,
  3.94,    3.94,    3.94,    3.94,
  3.37,    3.37,    3.37,    3.37,
  3.85,    3.85,    3.85,    3.85,
  3.52,    3.52,    3.52,    3.52,
  3.21,    3.21,    3.21,    3.21,
  3.39,    3.39,    3.39,    3.39,
  2.05,    2.05,    2.05,    2.05,
  2.59,    2.59,    2.59,    2.59,
  3.46,    3.46,    3.46,    3.46,
  3.07,    3.07,    3.07,    3.07,
  3.31,    3.31,    3.31,    3.31,
  3.53,    3.53,    3.53,    3.53,
  3.67,    3.67,    3.67,    3.67,
  3.76,    3.76,    3.76,    3.76,
  3.76,    3.76,    3.76,    3.76,
  3.67,    3.67,    3.67,    3.67,
  3.61,    3.61,    3.61,    3.61,
  3.58,    3.58,    3.58,    3.58,
  3.16,    3.16,    3.16,    3.16,
  3.32,    3.32,    3.32,    3.32,
  2.86,    2.86,    2.86,    2.86,
  2.39,    2.39,    2.39,    2.39,
  3.1,     3.1,     3.1,     3.1,
  2.82,    2.82,    2.82,    2.82,
  4.82,    4.82,    4.82,    4.82,
  4.74,    4.74,    4.74,    4.74,
  5.32,    5.32,    5.32,    5.32,
  4.68,    4.68,    4.68,    4.68,
  4.23,    4.23,    4.23,    4.23,
  3.95,    3.95,    3.95,    3.95,
  4.31,    4.31,    4.31,    4.31,
  4.2,     4.2,     4.2,     4.2,
  3.1,     3.1,     3.1,     3.1,
  2.56,    2.56,    2.56,    2.56,
  2.39,    2.39,    2.39,    2.39,
  2.07,    2.07,    2.07,    2.07,
  2.36,    2.36,    2.36,    2.36,
  1.97,    1.97,    1.97,    1.97,
  2.44,    2.44,    2.44,    2.44,
  2.26,    2.26,    2.26,    2.26,
  1.9,     1.9,     1.9,     1.9,
  2.14,    2.14,    2.14,    2.14,
  1.94,    1.94,    1.94,    1.94,
  0.78,    0.78,    0.78,    0.78,
  0.51,    0.51,    0.51,    0.51,
  1.39,    1.39,    1.39,    1.39,
  1.46,    1.46,    1.46,    1.46,
  1.53,    1.53,    1.53,    1.53,
  1.28,    1.28,    1.28,    1.28,
  1.01,    1.01,    1.01,    1.01,
  0.65,    0.65,    0.65,    0.65,
  0.94,    0.94,    0.94,    0.94,
  1.47,    1.47,    1.47,    1.47,
  1.11,    1.11,    1.11,    1.11,
  1.19,    1.19,    1.19,    1.19,
  0.87,    0.87,    0.87,    0.87,
  0.42,    0.42,    0.42,    0.42,
  0.54,    0.54,    0.54,    0.54,
  1.01,    1.01,    1.01,    1.01,
  0.97,    0.97,    0.97,    0.97,
  0.78,    0.78,    0.78,    0.78,
  1.23,    1.23,    1.23,    1.23,
  1.88,    1.88,    1.88,    1.88,
  2.04,    2.04,    2.04,    2.04,
  1.93,    1.93,    1.93,    1.93,
  2.03,    2.03,    2.03,    2.03,
  1.57,    1.57,    1.57,    1.57,
  1.57,    1.57,    1.57,    1.57,
  2.21,    2.21,    2.21,    2.21,
  2.64,    2.64,    2.64,    2.64,
  3.59,    3.59,    3.59,    3.59,
  3.46,    3.46,    3.46,    3.46,
  4.93,    4.93,    4.93,    4.93,
  3.67,    3.67,    3.67,    3.67,
  3.06,    3.06,    3.06,    3.06,
  4.11,    4.11,    4.11,    4.11,
  4.68,    4.68,    4.68,    4.68,
  4.91,    4.91,    4.91,    4.91,
  4.36,    4.36,    4.36,    4.36,
  4.37,    4.37,    4.37,    4.37,
  2.68,    2.68,    2.68,    2.68,
  2.98,    2.98,    2.98,    2.98,
  3.21,    3.21,    3.21,    3.21,
  2.9,     2.9,     2.9,     2.9,
  2.14,    2.14,    2.14,    2.14,
  2.5,     2.5,     2.5,     2.5,
  2.82,    2.82,    2.82,    2.82,
  1.75,    1.75,    1.75,    1.75,
  1.2,     1.2,     1.2,     1.2,
  1.05,    1.05,    1.05,    1.05,
  2.14,    2.14,    2.14,    2.14,
  2.41,    2.41,    2.41,    2.41,
  1.72,    1.72,    1.72,    1.72,
  1.96,    1.96,    1.96,    1.96,
  2.33,    2.33,    2.33,    2.33,
  1.92,    1.92,    1.92,    1.92,
  2.09,    2.09,    2.09,    2.09,
  2.39,    2.39,    2.39,    2.39,
  2.22,    2.22,    2.22,    2.22,
  2.38,    2.38,    2.38,    2.38,
  2.3,     2.3,     2.3,     2.3,
  2.47,    2.47,    2.47,    2.47,
  2.44,    2.44,    2.44,    2.44,
  2.22,    2.22,    2.22,    2.22,
  1.99,    1.99,    1.99,    1.99,
  1.58,    1.58,    1.58,    1.58,
  1.62,    1.62,    1.62,    1.62,
  1.82,    1.82,    1.82,    1.82,
  1.88,    1.88,    1.88,    1.88,
  2.17,    2.17,    2.17,    2.17,
  2.28,    2.28,    2.28,    2.28,
  2.81,    2.81,    2.81,    2.81,
  2.15,    2.15,    2.15,    2.15,
  2.69,    2.69,    2.69,    2.69,
  2.43,    2.43,    2.43,    2.43,
  2.78,    2.78,    2.78,    2.78,
  3.34,    3.34,    3.34,    3.34,
  3.39,    3.39,    3.39,    3.39,
  3.29,    3.29,    3.29,    3.29,
  3,       3,       3,       3,
  1.96,    1.96,    1.96,    1.96,
  1.97,    1.97,    1.97,    1.97,
  2.13,    2.13,    2.13,    2.13,
  1.44,    1.44,    1.44,    1.44,
  2.14,    2.14,    2.14,    2.14,
  2.87,    2.87,    2.87,    2.87,
  2.79,    2.79,    2.79,    2.79,
  1.78,    1.78,    1.78,    1.78,
  2.87,    2.87,    2.87,    2.87,
  3.39,    3.39,    3.39,    3.39,
  3.97,    3.97,    3.97,    3.97,
  3.21,    3.21,    3.21,    3.21,
  3.72,    3.72,    3.72,    3.72,
  2.99,    2.99,    2.99,    2.99,
  3.57,    3.57,    3.57,    3.57,
  2.3,     2.3,     2.3,     2.3,
  1.51,    1.51,    1.51,    1.51,
  0.86,    0.86,    0.86,    0.86,
  2.62,    2.62,    2.62,    2.62,
  1.63,    1.63,    1.63,    1.63,
  2.13,    2.13,    2.13,    2.13,
  1.42,    1.42,    1.42,    1.42,
  0.46,    0.46,    0.46,    0.46,
  1.59,    1.59,    1.59,    1.59,
  1.1,     1.1,     1.1,     1.1,
  1.4,     1.4,     1.4,     1.4,
  2.54,    2.54,    2.54,    2.54,
  2.04,    2.04,    2.04,    2.04,
  2.91,    2.91,    2.91,    2.91,
  2.5,     2.5,     2.5,     2.5,
  2.02,    2.02,    2.02,    2.02,
  2.14,    2.14,    2.14,    2.14,
  1.73,    1.73,    1.73,    1.73,
  1.84,    1.84,    1.84,    1.84,
  1.9,     1.9,     1.9,     1.9,
  2.42,    2.42,    2.42,    2.42,
  2.45,    2.45,    2.45,    2.45,
  2.51,    2.51,    2.51,    2.51,
  1.46,    1.46,    1.46,    1.46,
  2.04,    2.04,    2.04,    2.04,
  2.58,    2.58,    2.58,    2.58,
  3.31,    3.31,    3.31,    3.31,
  2.58,    2.58,    2.58,    2.58,
  1.81,    1.81,    1.81,    1.81,
  1.76,    1.76,    1.76,    1.76,
  2,       2,       2,       2,
  2.57,    2.57,    2.57,    2.57,
  1.97,    1.97,    1.97,    1.97,
  2.31,    2.31,    2.31,    2.31,
  3.1,     3.1,     3.1,     3.1,
  3.8,     3.8,     3.8,     3.8,
  4.17,    4.17,    4.17,    4.17,
  3.43,    3.43,    3.43,    3.43,
  2.98,    2.98,    2.98,    2.98,
  3.04,    3.04,    3.04,    3.04,
  2.27,    2.27,    2.27,    2.27,
  2.25,    2.25,    2.25,    2.25,
  2.67,    2.67,    2.67,    2.67,
  2.57,    2.57,    2.57,    2.57,
  2.51,    2.51,    2.51,    2.51,
  2.29,    2.29,    2.29,    2.29,
  1.85,    1.85,    1.85,    1.85,
  1.95,    1.95,    1.95,    1.95,
  2.22,    2.22,    2.22,    2.22,
  2.13,    2.13,    2.13,    2.13,
  1.92,    1.92,    1.92,    1.92,
  1.52,    1.52,    1.52,    1.52,
  1.63,    1.63,    1.63,    1.63,
  1.78,    1.78,    1.78,    1.78,
  1.92,    1.92,    1.92,    1.92,
  2.03,    2.03,    2.03,    2.03,
  1.86,    1.86,    1.86,    1.86,
  1.86,    1.86,    1.86,    1.86,
  2.05,    2.05,    2.05,    2.05,
  1.88,    1.88,    1.88,    1.88,
  2.14,    2.14,    2.14,    2.14,
  2.08,    2.08,    2.08,    2.08,
  1.88,    1.88,    1.88,    1.88,
  2.25,    2.25,    2.25,    2.25,
  2.38,    2.38,    2.38,    2.38,
  2.2,     2.2,     2.2,     2.2,
  2.12,    2.12,    2.12,    2.12,
  1.79,    1.79,    1.79,    1.79,
  2.13,    2.13,    2.13,    2.13,
  2.19,    2.19,    2.19,    2.19,
  2.74,    2.74,    2.74,    2.74,
  2.29,    2.29,    2.29,    2.29,
  2.22,    2.22,    2.22,    2.22,
  2.23,    2.23,    2.23,    2.23,
  2.1,     2.1,     2.1,     2.1,
  2.45,    2.45,    2.45,    2.45,
  2,       2,       2,       2,
  2.2,     2.2,     2.2,     2.2,
  1.63,    1.63,    1.63,    1.63,
  1.63,    1.63,    1.63,    1.63,
  1.97,    1.97,    1.97,    1.97,
  1.18,    1.18,    1.18,    1.18,
  1.28,    1.28,    1.28,    1.28,
  1.08,    1.08,    1.08,    1.08,
  0.71,    0.71,    0.71,    0.71,
  0.34,    0.34,    0.34,    0.34,
  0.64,    0.64,    0.64,    0.64,
  0.96,    0.96,    0.96,    0.96,
  0.63,    0.63,    0.63,    0.63,
  0.6,     0.6,     0.6,     0.6,
  1.18,    1.18,    1.18,    1.18,
  0.94,    0.94,    0.94,    0.94,
  1.39,    1.39,    1.39,    1.39,
  1.27,    1.27,    1.27,    1.27,
  0.88,    0.88,    0.88,    0.88,
  1.17,    1.17,    1.17,    1.17,
  1.4,     1.4,     1.4,     1.4,
  1.67,    1.67,    1.67,    1.67,
  2.06,    2.06,    2.06,    2.06,
  1.97,    1.97,    1.97,    1.97,
  1.49,    1.49,    1.49,    1.49,
  1.48,    1.48,    1.48,    1.48,
  1.32,    1.32,    1.32,    1.32,
  1.73,    1.73,    1.73,    1.73,
  1.51,    1.51,    1.51,    1.51,
  1.31,    1.31,    1.31,    1.31,
  1.2,     1.2,     1.2,     1.2,
  1.26,    1.26,    1.26,    1.26,
  1.57,    1.57,    1.57,    1.57,
  1.4,     1.4,     1.4,     1.4,
  1.69,    1.69,    1.69,    1.69,
  1.41,    1.41,    1.41,    1.41,
  1.02,    1.02,    1.02,    1.02,
  1.16,    1.16,    1.16,    1.16,
  1.93,    1.93,    1.93,    1.93,
  1.91,    1.91,    1.91,    1.91,
  1.57,    1.57,    1.57,    1.57,
  0.96,    0.96,    0.96,    0.96,
  1.46,    1.46,    1.46,    1.46,
  1.96,    1.96,    1.96,    1.96,
  1.98,    1.98,    1.98,    1.98,
  1.96,    1.96,    1.96,    1.96,
  2.18,    2.18,    2.18,    2.18,
  1.36,    1.36,    1.36,    1.36,
  1.26,    1.26,    1.26,    1.26,
  1.06,    1.06,    1.06,    1.06,
  1.07,    1.07,    1.07,    1.07,
  0.71,    0.71,    0.71,    0.71,
  1.3,     1.3,     1.3,     1.3,
  1.17,    1.17,    1.17,    1.17,
  2.31,    2.31,    2.31,    2.31,
  2.05,    2.05,    2.05,    2.05,
  2.02,    2.02,    2.02,    2.02,
  1.72,    1.72,    1.72,    1.72,
  1.72,    1.72,    1.72,    1.72,
  1.61,    1.61,    1.61,    1.61,
  1.71,    1.71,    1.71,    1.71,
  1.7,     1.7,     1.7,     1.7,
  1.72,    1.72,    1.72,    1.72,
  1.54,    1.54,    1.54,    1.54,
  1.29,    1.29,    1.29,    1.29,
  1.58,    1.58,    1.58,    1.58,
  1.57,    1.57,    1.57,    1.57,
  1.89,    1.89,    1.89,    1.89,
  1.81,    1.81,    1.81,    1.81,
  1.68,    1.68,    1.68,    1.68,
  1.71,    1.71,    1.71,    1.71,
  1.89,    1.89,    1.89,    1.89,
  2.05,    2.05,    2.05,    2.05,
  2.32,    2.32,    2.32,    2.32,
  2.28,    2.28,    2.28,    2.28,
  2.12,    2.12,    2.12,    2.12,
  2.19,    2.19,    2.19,    2.19,
  2.31,    2.31,    2.31,    2.31,
  2.34,    2.34,    2.34,    2.34,
  2.63,    2.63,    2.63,    2.63,
  2.4,     2.4,     2.4,     2.4,
  2.28,    2.28,    2.28,    2.28,
  2.29,    2.29,    2.29,    2.29,
  2.56,    2.56,    2.56,    2.56,
  2.47,    2.47,    2.47,    2.47,
  2.65,    2.65,    2.65,    2.65,
  2.55,    2.55,    2.55,    2.55,
  2.36,    2.36,    2.36,    2.36,
  2.76,    2.76,    2.76,    2.76,
  2.6,     2.6,     2.6,     2.6,
  2.77,    2.77,    2.77,    2.77,
  2.44,    2.44,    2.44,    2.44,
  1.92,    1.92,    1.92,    1.92,
  2.42,    2.42,    2.42,    2.42,
  1.82,    1.82,    1.82,    1.82,
  2.01,    2.01,    2.01,    2.01,
  2.36,    2.36,    2.36,    2.36,
  2.3,     2.3,     2.3,     2.3,
  2.34,    2.34,    2.34,    2.34,
  2.29,    2.29,    2.29,    2.29,
  1.9,     1.9,     1.9,     1.9,
  2.5,     2.5,     2.5,     2.5,
  2.53,    2.53,    2.53,    2.53,
  2.48,    2.48,    2.48,    2.48,
  2.95,    2.95,    2.95,    2.95,
  2.78,    2.78,    2.78,    2.78,
  2.48,    2.48,    2.48,    2.48,
  3.04,    3.04,    3.04,    3.04,
  2.1,     2.1,     2.1,     2.1,
  2.14,    2.14,    2.14,    2.14,
  1.86,    1.86,    1.86,    1.86,
  2.19,    2.19,    2.19,    2.19,
  2.18,    2.18,    2.18,    2.18,
  2.06,    2.06,    2.06,    2.06,
  1.78,    1.78,    1.78,    1.78,
  1.97,    1.97,    1.97,    1.97,
  2.19,    2.19,    2.19,    2.19,
  2.36,    2.36,    2.36,    2.36,
  2.52,    2.52,    2.52,    2.52,
  2.17,    2.17,    2.17,    2.17,
  2.16,    2.16,    2.16,    2.16,
  2.18,    2.18,    2.18,    2.18,
  1.9,     1.9,     1.9,     1.9,
  2.33,    2.33,    2.33,    2.33,
  2.52,    2.52,    2.52,    2.52,
  2.5,     2.5,     2.5,     2.5,
  2.39,    2.39,    2.39,    2.39,
  2.65,    2.65,    2.65,    2.65,
  2.64,    2.64,    2.64,    2.64,
  2.82,    2.82,    2.82,    2.82,
  2.5,     2.5,     2.5,     2.5,
  2.39,    2.39,    2.39,    2.39,
  2.5,     2.5,     2.5,     2.5,
  2.34,    2.34,    2.34,    2.34,
  2.2,     2.2,     2.2,     2.2,
  2.04,    2.04,    2.04,    2.04,
  2.46,    2.46,    2.46,    2.46,
  2.19,    2.19,    2.19,    2.19,
  2.34,    2.34,    2.34,    2.34,
  2.55,    2.55,    2.55,    2.55,
  2.76,    2.76,    2.76,    2.76,
  3.17,    3.17,    3.17,    3.17,
  2.46,    2.46,    2.46,    2.46,
  2.52,    2.52,    2.52,    2.52,
  2.74,    2.74,    2.74,    2.74,
  2.8,     2.8,     2.8,     2.8,
  2.68,    2.68,    2.68,    2.68,
  3.23,    3.23,    3.23,    3.23,
  3.19,    3.19,    3.19,    3.19,
  2.64,    2.64,    2.64,    2.64,
  2.82,    2.82,    2.82,    2.82,
  2.64,    2.64,    2.64,    2.64,
  2.82,    2.82,    2.82,    2.82,
  2.67,    2.67,    2.67,    2.67,
  2.89,    2.89,    2.89,    2.89,
  2.25,    2.25,    2.25,    2.25,
  3.07,    3.07,    3.07,    3.07,
  2.75,    2.75,    2.75,    2.75,
  2.55,    2.55,    2.55,    2.55,
  2.49,    2.49,    2.49,    2.49,
  1.62,    1.62,    1.62,    1.62,
  1.89,    1.89,    1.89,    1.89,
  2.29,    2.29,    2.29,    2.29,
  2.54,    2.54,    2.54,    2.54,
  2.03,    2.03,    2.03,    2.03,
  1.97,    1.97,    1.97,    1.97,
  1.88,    1.88,    1.88,    1.88,
  1.81,    1.81,    1.81,    1.81,
  1.96,    1.96,    1.96,    1.96,
  2.32,    2.32,    2.32,    2.32,
  2.03,    2.03,    2.03,    2.03,
  2.06,    2.06,    2.06,    2.06,
  1.99,    1.99,    1.99,    1.99,
  1.86,    1.86,    1.86,    1.86,
  2.12,    2.12,    2.12,    2.12,
  1.98,    1.98,    1.98,    1.98,
  1.81,    1.81,    1.81,    1.81,
  1.66,    1.66,    1.66,    1.66,
  1.76,    1.76,    1.76,    1.76,
  2.23,    2.23,    2.23,    2.23,
  2.13,    2.13,    2.13,    2.13,
  1.78,    1.78,    1.78,    1.78,
  1.61,    1.61,    1.61,    1.61,
  1.52,    1.52,    1.52,    1.52,
  1.98,    1.98,    1.98,    1.98,
  2.07,    2.07,    2.07,    2.07,
  2.15,    2.15,    2.15,    2.15,
  2.36,    2.36,    2.36,    2.36,
  2.23,    2.23,    2.23,    2.23,
  2,       2,       2,       2,
  1.93,    1.93,    1.93,    1.93,
  1.96,    1.96,    1.96,    1.96,
  1.79,    1.79,    1.79,    1.79,
  1.34,    1.34,    1.34,    1.34,
  1.81,    1.81,    1.81,    1.81,
  1.5,     1.5,     1.5,     1.5,
  1.25,    1.25,    1.25,    1.25,
  1.52,    1.52,    1.52,    1.52,
  1.32,    1.32,    1.32,    1.32,
  1.56,    1.56,    1.56,    1.56,
  1.65,    1.65,    1.65,    1.65,
  1.37,    1.37,    1.37,    1.37,
  1.21,    1.21,    1.21,    1.21,
  1.62,    1.62,    1.62,    1.62,
  1.27,    1.27,    1.27,    1.27,
  0.98,    0.98,    0.98,    0.98,
  0.88,    0.88,    0.88,    0.88,
  1.09,    1.09,    1.09,    1.09,
  0.95,    0.95,    0.95,    0.95,
  1.13,    1.13,    1.13,    1.13,
  1.48,    1.48,    1.48,    1.48,
  0.27,    0.27,    0.27,    0.27,
  0.62,    0.62,    0.62,    0.62,
  1.5,     1.5,     1.5,     1.5,
  1.66,    1.66,    1.66,    1.66,
  1.65,    1.65,    1.65,    1.65,
  1.74,    1.74,    1.74,    1.74,
  1.37,    1.37,    1.37,    1.37,
  1.26,    1.26,    1.26,    1.26,
  1.38,    1.38,    1.38,    1.38,
  1.11,    1.11,    1.11,    1.11,
  1.22,    1.22,    1.22,    1.22,
  1.85,    1.85,    1.85,    1.85,
  2.31,    2.31,    2.31,    2.31,
  1.74,    1.74,    1.74,    1.74,
  2.02,    2.02,    2.02,    2.02,
  2.08,    2.08,    2.08,    2.08,
  2.4,     2.4,     2.4,     2.4,
  2.77,    2.77,    2.77,    2.77,
  2.69,    2.69,    2.69,    2.69,
  2.79,    2.79,    2.79,    2.79,
  2.8,     2.8,     2.8,     2.8,
  2.64,    2.64,    2.64,    2.64,
  2.73,    2.73,    2.73,    2.73,
  3.06,    3.06,    3.06,    3.06,
  3.93,    3.93,    3.93,    3.93,
  3.63,    3.63,    3.63,    3.63,
  3.07,    3.07,    3.07,    3.07,
  3.74,    3.74,    3.74,    3.74,
  5.02,    5.02,    5.02,    5.02,
  4.14,    4.14,    4.14,    4.14,
  4.3,     4.3,     4.3,     4.3,
  4.57,    4.57,    4.57,    4.57,
  4.57,    4.57,    4.57,    4.57,
  3.68,    3.68,    3.68,    3.68,
  4.36,    4.36,    4.36,    4.36,
  4.14,    4.14,    4.14,    4.14,
  4.55,    4.55,    4.55,    4.55,
  4.06,    4.06,    4.06,    4.06,
  4.23,    4.23,    4.23,    4.23,
  3.89,    3.89,    3.89,    3.89,
  4.21,    4.21,    4.21,    4.21,
  3.7,     3.7,     3.7,     3.7,
  3.9,     3.9,     3.9,     3.9,
  3.76,    3.76,    3.76,    3.76,
  3.05,    3.05,    3.05,    3.05,
  3.11,    3.11,    3.11,    3.11,
  2.44,    2.44,    2.44,    2.44,
  2.21,    2.21,    2.21,    2.21,
  2.01,    2.01,    2.01,    2.01,
  2.29,    2.29,    2.29,    2.29,
  2.11,    2.11,    2.11,    2.11,
  2.62,    2.62,    2.62,    2.62,
  2.46,    2.46,    2.46,    2.46,
  2.52,    2.52,    2.52,    2.52,
  2.04,    2.04,    2.04,    2.04,
  2.45,    2.45,    2.45,    2.45,
  2.86,    2.86,    2.86,    2.86,
  2.76,    2.76,    2.76,    2.76,
  2.56,    2.56,    2.56,    2.56,
  2.66,    2.66,    2.66,    2.66,
  2.66,    2.66,    2.66,    2.66,
  2.66,    2.66,    2.66,    2.66,
  2.78,    2.78,    2.78,    2.78,
  2.82,    2.82,    2.82,    2.82,
  2.94,    2.94,    2.94,    2.94,
  2.91,    2.91,    2.91,    2.91,
  2.63,    2.63,    2.63,    2.63,
  2.72,    2.72,    2.72,    2.72,
  2.64,    2.64,    2.64,    2.64,
  2.49,    2.49,    2.49,    2.49,
  2.68,    2.68,    2.68,    2.68,
  2.83,    2.83,    2.83,    2.83,
  3,       3,       3,       3,
  3.03,    3.03,    3.03,    3.03,
  2.67,    2.67,    2.67,    2.67,
  2.66,    2.66,    2.66,    2.66,
  2.67,    2.67,    2.67,    2.67,
  2.71,    2.71,    2.71,    2.71,
  2.96,    2.96,    2.96,    2.96,
  2.77,    2.77,    2.77,    2.77,
  3.46,    3.46,    3.46,    3.46,
  2.88,    2.88,    2.88,    2.88,
  3.44,    3.44,    3.44,    3.44,
  3.53,    3.53,    3.53,    3.53,
  3.78,    3.78,    3.78,    3.78,
  4.03,    4.03,    4.03,    4.03,
  3.69,    3.69,    3.69,    3.69,
  3.53,    3.53,    3.53,    3.53,
  3.48,    3.48,    3.48,    3.48,
  3.83,    3.83,    3.83,    3.83,
  3.43,    3.43,    3.43,    3.43,
  3.64,    3.64,    3.64,    3.64,
  2.59,    2.59,    2.59,    2.59,
  2.3,     2.3,     2.3,     2.3,
  2.05,    2.05,    2.05,    2.05,
  1.99,    1.99,    1.99,    1.99,
  2.17,    2.17,    2.17,    2.17,
  2.27,    2.27,    2.27,    2.27,
  2.31,    2.31,    2.31,    2.31,
  2.9,     2.9,     2.9,     2.9,
  3.1,     3.1,     3.1,     3.1,
  2.59,    2.59,    2.59,    2.59,
  3.13,    3.13,    3.13,    3.13,
  3.04,    3.04,    3.04,    3.04,
  3.11,    3.11,    3.11,    3.11,
  3.25,    3.25,    3.25,    3.25,
  3.04,    3.04,    3.04,    3.04,
  2.78,    2.78,    2.78,    2.78,
  2.05,    2.05,    2.05,    2.05,
  2.04,    2.04,    2.04,    2.04,
  2.44,    2.44,    2.44,    2.44,
  2.4,     2.4,     2.4,     2.4,
  2.67,    2.67,    2.67,    2.67,
  2.67,    2.67,    2.67,    2.67,
  2.3,     2.3,     2.3,     2.3,
  2.49,    2.49,    2.49,    2.49,
  2.9,     2.9,     2.9,     2.9,
  2.86,    2.86,    2.86,    2.86,
  2.48,    2.48,    2.48,    2.48,
  2.39,    2.39,    2.39,    2.39,
  2.44,    2.44,    2.44,    2.44,
  2.34,    2.34,    2.34,    2.34,
  1.95,    1.95,    1.95,    1.95,
  1.98,    1.98,    1.98,    1.98,
  1.8,     1.8,     1.8,     1.8,
  1.77,    1.77,    1.77,    1.77,
  1.71,    1.71,    1.71,    1.71,
  1.35,    1.35,    1.35,    1.35,
  0.87,    0.87,    0.87,    0.87,
  0.5,     0.5,     0.5,     0.5,
  1.06,    1.06,    1.06,    1.06,
  1.04,    1.04,    1.04,    1.04,
  1.75,    1.75,    1.75,    1.75,
  1.69,    1.69,    1.69,    1.69,
  1.54,    1.54,    1.54,    1.54,
  1.42,    1.42,    1.42,    1.42,
  1.13,    1.13,    1.13,    1.13,
  0.73,    0.73,    0.73,    0.73,
  1.03,    1.03,    1.03,    1.03,
  1.04,    1.04,    1.04,    1.04,
  1.43,    1.43,    1.43,    1.43,
  1.55,    1.55,    1.55,    1.55,
  2.2,     2.2,     2.2,     2.2,
  2.06,    2.06,    2.06,    2.06,
  1.45,    1.45,    1.45,    1.45,
  1.45,    1.45,    1.45,    1.45,
  1.44,    1.44,    1.44,    1.44,
  1.51,    1.51,    1.51,    1.51,
  0.47,    0.47,    0.47,    0.47,
  0.34,    0.34,    0.34,    0.34,
  0.83,    0.83,    0.83,    0.83,
  0.51,    0.51,    0.51,    0.51,
  1.41,    1.41,    1.41,    1.41,
  0.54,    0.54,    0.54,    0.54,
  0.29,    0.29,    0.29,    0.29,
  0.62,    0.62,    0.62,    0.62,
  0.38,    0.38,    0.38,    0.38,
  1.18,    1.18,    1.18,    1.18,
  1.18,    1.18,    1.18,    1.18,
  1.03,    1.03,    1.03,    1.03,
  1.08,    1.08,    1.08,    1.08,
  1.98,    1.98,    1.98,    1.98,
  1.05,    1.05,    1.05,    1.05,
  0.83,    0.83,    0.83,    0.83,
  1.01,    1.01,    1.01,    1.01,
  1,       1,       1,       1,
  1.01,    1.01,    1.01,    1.01,
  1.38,    1.38,    1.38,    1.38,
  0.3,     0.3,     0.3,     0.3,
  0.66,    0.66,    0.66,    0.66,
  0.61,    0.61,    0.61,    0.61,
  0.57,    0.57,    0.57,    0.57,
  0.81,    0.81,    0.81,    0.81,
  0.8,     0.8,     0.8,     0.8,
  0.54,    0.54,    0.54,    0.54,
  0.7,     0.7,     0.7,     0.7,
  0.69,    0.69,    0.69,    0.69,
  0.63,    0.63,    0.63,    0.63,
  0.78,    0.78,    0.78,    0.78,
  1.84,    1.84,    1.84,    1.84,
  2.54,    2.54,    2.54,    2.54,
  2.23,    2.23,    2.23,    2.23,
  1.71,    1.71,    1.71,    1.71,
  3.62,    3.62,    3.62,    3.62,
  2.49,    2.49,    2.49,    2.49,
  2.27,    2.27,    2.27,    2.27,
  2.22,    2.22,    2.22,    2.22,
  2.16,    2.16,    2.16,    2.16,
  2.1,     2.1,     2.1,     2.1,
  1.81,    1.81,    1.81,    1.81,
  1.73,    1.73,    1.73,    1.73,
  2.02,    2.02,    2.02,    2.02,
  2.02,    2.02,    2.02,    2.02,
  1.99,    1.99,    1.99,    1.99,
  1.54,    1.54,    1.54,    1.54,
  1.7,     1.7,     1.7,     1.7,
  1.48,    1.48,    1.48,    1.48,
  1.61,    1.61,    1.61,    1.61,
  1.86,    1.86,    1.86,    1.86,
  2.04,    2.04,    2.04,    2.04,
  1.77,    1.77,    1.77,    1.77,
  1.92,    1.92,    1.92,    1.92,
  2.12,    2.12,    2.12,    2.12,
  1.64,    1.64,    1.64,    1.64,
  1.82,    1.82,    1.82,    1.82,
  2.02,    2.02,    2.02,    2.02,
  1.87,    1.87,    1.87,    1.87,
  1.73,    1.73,    1.73,    1.73,
  1.99,    1.99,    1.99,    1.99,
  1.89,    1.89,    1.89,    1.89,
  1.68,    1.68,    1.68,    1.68,
  1.36,    1.36,    1.36,    1.36,
  1.96,    1.96,    1.96,    1.96,
  1.93,    1.93,    1.93,    1.93,
  1.59,    1.59,    1.59,    1.59,
  1.18,    1.18,    1.18,    1.18,
  1.35,    1.35,    1.35,    1.35,
  1.59,    1.59,    1.59,    1.59,
  2.24,    2.24,    2.24,    2.24,
  1.98,    1.98,    1.98,    1.98,
  1.61,    1.61,    1.61,    1.61,
  1.25,    1.25,    1.25,    1.25,
  1.7,     1.7,     1.7,     1.7,
  1.86,    1.86,    1.86,    1.86,
  0.89,    0.89,    0.89,    0.89,
  0.96,    0.96,    0.96,    0.96,
  1.56,    1.56,    1.56,    1.56,
  2.63,    2.63,    2.63,    2.63,
  2.69,    2.69,    2.69,    2.69,
  2.73,    2.73,    2.73,    2.73,
  3.74,    3.74,    3.74,    3.74,
  2.35,    2.35,    2.35,    2.35,
  3.03,    3.03,    3.03,    3.03,
  3.13,    3.13,    3.13,    3.13,
  2.86,    2.86,    2.86,    2.86,
  2.59,    2.59,    2.59,    2.59,
  2.25,    2.25,    2.25,    2.25,
  2.11,    2.11,    2.11,    2.11,
  1.96,    1.96,    1.96,    1.96,
  1.81,    1.81,    1.81,    1.81,
  1.54,    1.54,    1.54,    1.54,
  1.85,    1.85,    1.85,    1.85,
  1.81,    1.81,    1.81,    1.81,
  1.93,    1.93,    1.93,    1.93,
  1.88,    1.88,    1.88,    1.88,
  1.88,    1.88,    1.88,    1.88,
  1.92,    1.92,    1.92,    1.92,
  1.85,    1.85,    1.85,    1.85,
  1.82,    1.82,    1.82,    1.82,
  1.85,    1.85,    1.85,    1.85,
  1.76,    1.76,    1.76,    1.76,
  1.63,    1.63,    1.63,    1.63,
  1.72,    1.72,    1.72,    1.72,
  1.89,    1.89,    1.89,    1.89,
  2.1,     2.1,     2.1,     2.1,
  2.22,    2.22,    2.22,    2.22,
  2.01,    2.01,    2.01,    2.01,
  2.02,    2.02,    2.02,    2.02,
  2.2,     2.2,     2.2,     2.2,
  2.31,    2.31,    2.31,    2.31,
  1.92,    1.92,    1.92,    1.92,
  2.31,    2.31,    2.31,    2.31,
  2.29,    2.29,    2.29,    2.29,
  2.06,    2.06,    2.06,    2.06,
  2.16,    2.16,    2.16,    2.16,
  2.1,     2.1,     2.1,     2.1,
  1.95,    1.95,    1.95,    1.95,
  2.47,    2.47,    2.47,    2.47,
  2.45,    2.45,    2.45,    2.45,
  2.28,    2.28,    2.28,    2.28,
  2.5,     2.5,     2.5,     2.5,
  2.55,    2.55,    2.55,    2.55,
  2.52,    2.52,    2.52,    2.52,
  2.66,    2.66,    2.66,    2.66,
  3.07,    3.07,    3.07,    3.07,
  2.86,    2.86,    2.86,    2.86,
  3.25,    3.25,    3.25,    3.25,
  4.26,    4.26,    4.26,    4.26,
  4.44,    4.44,    4.44,    4.44,
  4.33,    4.33,    4.33,    4.33,
  4.13,    4.13,    4.13,    4.13,
  3.21,    3.21,    3.21,    3.21,
  3.66,    3.66,    3.66,    3.66,
  3.79,    3.79,    3.79,    3.79,
  3.42,    3.42,    3.42,    3.42,
  2.93,    2.93,    2.93,    2.93,
  1.79,    1.79,    1.79,    1.79,
  1.49,    1.49,    1.49,    1.49,
  1.5,     1.5,     1.5,     1.5,
  1.3,     1.3,     1.3,     1.3,
  1.01,    1.01,    1.01,    1.01,
  1.11,    1.11,    1.11,    1.11,
  1.21,    1.21,    1.21,    1.21,
  1.07,    1.07,    1.07,    1.07,
  1.26,    1.26,    1.26,    1.26,
  1.06,    1.06,    1.06,    1.06,
  0.97,    0.97,    0.97,    0.97,
  0.86,    0.86,    0.86,    0.86,
  1.22,    1.22,    1.22,    1.22,
  1.4,     1.4,     1.4,     1.4,
  1.55,    1.55,    1.55,    1.55,
  1.63,    1.63,    1.63,    1.63,
  1.59,    1.59,    1.59,    1.59,
  1.27,    1.27,    1.27,    1.27,
  1.15,    1.15,    1.15,    1.15,
  0.51,    0.51,    0.51,    0.51,
  1.51,    1.51,    1.51,    1.51,
  1.5,     1.5,     1.5,     1.5,
  1.62,    1.62,    1.62,    1.62,
  0.91,    0.91,    0.91,    0.91,
  1.14,    1.14,    1.14,    1.14,
  0.95,    0.95,    0.95,    0.95,
  1.15,    1.15,    1.15,    1.15,
  1.24,    1.24,    1.24,    1.24,
  1.3,     1.3,     1.3,     1.3,
  1.35,    1.35,    1.35,    1.35,
  0.4,     0.4,     0.4,     0.4,
  1.01,    1.01,    1.01,    1.01,
  1.62,    1.62,    1.62,    1.62,
  1.89,    1.89,    1.89,    1.89,
  1.71,    1.71,    1.71,    1.71,
  2.52,    2.52,    2.52,    2.52,
  2.4,     2.4,     2.4,     2.4,
  2.32,    2.32,    2.32,    2.32,
  2.58,    2.58,    2.58,    2.58,
  2.47,    2.47,    2.47,    2.47,
  3.18,    3.18,    3.18,    3.18,
  2.43,    2.43,    2.43,    2.43,
  2.04,    2.04,    2.04,    2.04,
  1.69,    1.69,    1.69,    1.69,
  1.79,    1.79,    1.79,    1.79,
  1.47,    1.47,    1.47,    1.47,
  0.86,    0.86,    0.86,    0.86,
  0.73,    0.73,    0.73,    0.73,
  0.31,    0.31,    0.31,    0.31,
  0.46,    0.46,    0.46,    0.46,
  0.96,    0.96,    0.96,    0.96,
  1.19,    1.19,    1.19,    1.19,
  1.19,    1.19,    1.19,    1.19,
  1.27,    1.27,    1.27,    1.27,
  1.1,     1.1,     1.1,     1.1,
  0.97,    0.97,    0.97,    0.97,
  1.2,     1.2,     1.2,     1.2,
  1.3,     1.3,     1.3,     1.3,
  1.24,    1.24,    1.24,    1.24,
  1.27,    1.27,    1.27,    1.27,
  1.46,    1.46,    1.46,    1.46,
  1.79,    1.79,    1.79,    1.79,
  1.65,    1.65,    1.65,    1.65,
  2.04,    2.04,    2.04,    2.04,
  2.16,    2.16,    2.16,    2.16,
  1.99,    1.99,    1.99,    1.99,
  2.13,    2.13,    2.13,    2.13,
  2.41,    2.41,    2.41,    2.41,
  2.15,    2.15,    2.15,    2.15,
  2.46,    2.46,    2.46,    2.46,
  2.56,    2.56,    2.56,    2.56,
  3.16,    3.16,    3.16,    3.16,
  2.54,    2.54,    2.54,    2.54,
  2.4,     2.4,     2.4,     2.4,
  2.55,    2.55,    2.55,    2.55,
  2.73,    2.73,    2.73,    2.73,
  2.64,    2.64,    2.64,    2.64,
  2.41,    2.41,    2.41,    2.41,
  2.51,    2.51,    2.51,    2.51,
  2.5,     2.5,     2.5,     2.5,
  2.31,    2.31,    2.31,    2.31,
  3.33,    3.33,    3.33,    3.33,
  3.58,    3.58,    3.58,    3.58,
  3.89,    3.89,    3.89,    3.89,
  4.05,    4.05,    4.05,    4.05,
  4.54,    4.54,    4.54,    4.54,
  4.37,    4.37,    4.37,    4.37,
  4.12,    4.12,    4.12,    4.12,
  4.01,    4.01,    4.01,    4.01,
  4.68,    4.68,    4.68,    4.68,
  4.33,    4.33,    4.33,    4.33,
  4.21,    4.21,    4.21,    4.21,
  4.1,     4.1,     4.1,     4.1,
  4.07,    4.07,    4.07,    4.07,
  3.5,     3.5,     3.5,     3.5,
  2.74,    2.74,    2.74,    2.74,
  2.53,    2.53,    2.53,    2.53,
  2.48,    2.48,    2.48,    2.48,
  2.88,    2.88,    2.88,    2.88,
  2.88,    2.88,    2.88,    2.88,
  3,       3,       3,       3,
  3.15,    3.15,    3.15,    3.15,
  3.03,    3.03,    3.03,    3.03,
  3.07,    3.07,    3.07,    3.07,
  3.1,     3.1,     3.1,     3.1,
  3.04,    3.04,    3.04,    3.04,
  3.01,    3.01,    3.01,    3.01,
  2.88,    2.88,    2.88,    2.88,
  2.83,    2.83,    2.83,    2.83,
  2.75,    2.75,    2.75,    2.75,
  2.72,    2.72,    2.72,    2.72,
  2.65,    2.65,    2.65,    2.65,
  2.8,     2.8,     2.8,     2.8,
  2.67,    2.67,    2.67,    2.67,
  2.65,    2.65,    2.65,    2.65,
  2.29,    2.29,    2.29,    2.29,
  2.32,    2.32,    2.32,    2.32,
  2.6,     2.6,     2.6,     2.6,
  2.72,    2.72,    2.72,    2.72,
  2.58,    2.58,    2.58,    2.58,
  1.54,    1.54,    1.54,    1.54,
  1.36,    1.36,    1.36,    1.36,
  2.12,    2.12,    2.12,    2.12,
  2.16,    2.16,    2.16,    2.16,
  2.21,    2.21,    2.21,    2.21,
  1.86,    1.86,    1.86,    1.86,
  2.16,    2.16,    2.16,    2.16,
  1.4,     1.4,     1.4,     1.4,
  1.42,    1.42,    1.42,    1.42,
  2.36,    2.36,    2.36,    2.36,
  2.19,    2.19,    2.19,    2.19,
  3.09,    3.09,    3.09,    3.09,
  3.7,     3.7,     3.7,     3.7,
  3.78,    3.78,    3.78,    3.78,
  3.99,    3.99,    3.99,    3.99,
  3.62,    3.62,    3.62,    3.62,
  3.92,    3.92,    3.92,    3.92,
  3.54,    3.54,    3.54,    3.54,
  3.58,    3.58,    3.58,    3.58,
  3.34,    3.34,    3.34,    3.34,
  3.24,    3.24,    3.24,    3.24,
  3.16,    3.16,    3.16,    3.16,
  2.89,    2.89,    2.89,    2.89,
  2.37,    2.37,    2.37,    2.37,
  2.54,    2.54,    2.54,    2.54,
  2.79,    2.79,    2.79,    2.79,
  2.63,    2.63,    2.63,    2.63,
  2.82,    2.82,    2.82,    2.82,
  3.05,    3.05,    3.05,    3.05,
  2.92,    2.92,    2.92,    2.92,
  2.52,    2.52,    2.52,    2.52,
  2.05,    2.05,    2.05,    2.05,
  2.13,    2.13,    2.13,    2.13,
  2.59,    2.59,    2.59,    2.59,
  3.13,    3.13,    3.13,    3.13,
  2.86,    2.86,    2.86,    2.86,
  2.82,    2.82,    2.82,    2.82,
  2.52,    2.52,    2.52,    2.52,
  2.52,    2.52,    2.52,    2.52,
  2.33,    2.33,    2.33,    2.33,
  2.92,    2.92,    2.92,    2.92,
  2.29,    2.29,    2.29,    2.29,
  2.64,    2.64,    2.64,    2.64,
  2.46,    2.46,    2.46,    2.46,
  2.74,    2.74,    2.74,    2.74,
  1.18,    1.18,    1.18,    1.18,
  2.07,    2.07,    2.07,    2.07,
  2.37,    2.37,    2.37,    2.37,
  2.44,    2.44,    2.44,    2.44,
  2.28,    2.28,    2.28,    2.28,
  2.57,    2.57,    2.57,    2.57,
  2.2,     2.2,     2.2,     2.2,
  1.95,    1.95,    1.95,    1.95,
  2.32,    2.32,    2.32,    2.32,
  1.97,    1.97,    1.97,    1.97,
  1.47,    1.47,    1.47,    1.47,
  0.8,     0.8,     0.8,     0.8,
  1,       1,       1,       1,
  1.18,    1.18,    1.18,    1.18,
  1.34,    1.34,    1.34,    1.34,
  1.33,    1.33,    1.33,    1.33,
  1.33,    1.33,    1.33,    1.33,
  1.53,    1.53,    1.53,    1.53,
  1.77,    1.77,    1.77,    1.77,
  1.24,    1.24,    1.24,    1.24,
  0.8,     0.8,     0.8,     0.8,
  0.78,    0.78,    0.78,    0.78,
  0.88,    0.88,    0.88,    0.88,
  1.24,    1.24,    1.24,    1.24,
  0.8,     0.8,     0.8,     0.8,
  1.98,    1.98,    1.98,    1.98,
  2.29,    2.29,    2.29,    2.29,
  2.37,    2.37,    2.37,    2.37,
  2.38,    2.38,    2.38,    2.38,
  2.29,    2.29,    2.29,    2.29,
  2.64,    2.64,    2.64,    2.64,
  2.7,     2.7,     2.7,     2.7,
  2.59,    2.59,    2.59,    2.59,
  2.55,    2.55,    2.55,    2.55,
  2.4,     2.4,     2.4,     2.4,
  2.49,    2.49,    2.49,    2.49,
  2.2,     2.2,     2.2,     2.2,
  1.95,    1.95,    1.95,    1.95,
  2.19,    2.19,    2.19,    2.19,
  1.96,    1.96,    1.96,    1.96,
  2.31,    2.31,    2.31,    2.31,
  2.64,    2.64,    2.64,    2.64,
  2.4,     2.4,     2.4,     2.4,
  2.58,    2.58,    2.58,    2.58,
  2.37,    2.37,    2.37,    2.37,
  2.39,    2.39,    2.39,    2.39,
  2.13,    2.13,    2.13,    2.13,
  1.75,    1.75,    1.75,    1.75,
  1.88,    1.88,    1.88,    1.88,
  2.65,    2.65,    2.65,    2.65,
  1.89,    1.89,    1.89,    1.89,
  2.06,    2.06,    2.06,    2.06,
  1.81,    1.81,    1.81,    1.81,
  2.06,    2.06,    2.06,    2.06,
  1.97,    1.97,    1.97,    1.97,
  1.76,    1.76,    1.76,    1.76,
  1.65,    1.65,    1.65,    1.65,
  1.64,    1.64,    1.64,    1.64,
  1.46,    1.46,    1.46,    1.46,
  1.03,    1.03,    1.03,    1.03,
  1.49,    1.49,    1.49,    1.49,
  1.22,    1.22,    1.22,    1.22,
  0.75,    0.75,    0.75,    0.75,
  0.53,    0.53,    0.53,    0.53,
  0.58,    0.58,    0.58,    0.58,
  0.59,    0.59,    0.59,    0.59,
  0.55,    0.55,    0.55,    0.55,
  0.53,    0.53,    0.53,    0.53,
  0.64,    0.64,    0.64,    0.64,
  0.34,    0.34,    0.34,    0.34,
  0.67,    0.67,    0.67,    0.67,
  0.91,    0.91,    0.91,    0.91,
  1.83,    1.83,    1.83,    1.83,
  1.89,    1.89,    1.89,    1.89,
  2.27,    2.27,    2.27,    2.27,
  2.1,     2.1,     2.1,     2.1,
  2.17,    2.17,    2.17,    2.17,
  2.37,    2.37,    2.37,    2.37,
  2.42,    2.42,    2.42,    2.42,
  3.05,    3.05,    3.05,    3.05,
  2.87,    2.87,    2.87,    2.87,
  3.03,    3.03,    3.03,    3.03,
  2.78,    2.78,    2.78,    2.78,
  3.25,    3.25,    3.25,    3.25,
  3.51,    3.51,    3.51,    3.51,
  3.28,    3.28,    3.28,    3.28,
  3.4,     3.4,     3.4,     3.4,
  3.45,    3.45,    3.45,    3.45,
  3.47,    3.47,    3.47,    3.47,
  3.33,    3.33,    3.33,    3.33,
  3.32,    3.32,    3.32,    3.32,
  3.4,     3.4,     3.4,     3.4,
  2.91,    2.91,    2.91,    2.91,
  2.71,    2.71,    2.71,    2.71,
  3.1,     3.1,     3.1,     3.1,
  2.84,    2.84,    2.84,    2.84,
  2.61,    2.61,    2.61,    2.61,
  2.4,     2.4,     2.4,     2.4,
  2.23,    2.23,    2.23,    2.23,
  2.23,    2.23,    2.23,    2.23,
  2.5,     2.5,     2.5,     2.5,
  2.82,    2.82,    2.82,    2.82,
  2.99,    2.99,    2.99,    2.99,
  2.96,    2.96,    2.96,    2.96,
  2.95,    2.95,    2.95,    2.95,
  2.87,    2.87,    2.87,    2.87,
  2.86,    2.86,    2.86,    2.86,
  3.03,    3.03,    3.03,    3.03,
  3.71,    3.71,    3.71,    3.71,
  3.18,    3.18,    3.18,    3.18,
  3.9,     3.9,     3.9,     3.9,
  4.33,    4.33,    4.33,    4.33,
  3.98,    3.98,    3.98,    3.98,
  3.68,    3.68,    3.68,    3.68,
  3.35,    3.35,    3.35,    3.35,
  3.1,     3.1,     3.1,     3.1,
  3.4,     3.4,     3.4,     3.4,
  3.97,    3.97,    3.97,    3.97,
  3.5,     3.5,     3.5,     3.5,
  3.32,    3.32,    3.32,    3.32,
  3.41,    3.41,    3.41,    3.41,
  3.29,    3.29,    3.29,    3.29,
  2.9,     2.9,     2.9,     2.9,
  2.66,    2.66,    2.66,    2.66,
  2.59,    2.59,    2.59,    2.59,
  2.91,    2.91,    2.91,    2.91,
  2.42,    2.42,    2.42,    2.42,
  1.88,    1.88,    1.88,    1.88,
  2.74,    2.74,    2.74,    2.74,
  2.61,    2.61,    2.61,    2.61,
  2.58,    2.58,    2.58,    2.58,
  2.15,    2.15,    2.15,    2.15,
  2.26,    2.26,    2.26,    2.26,
  2.65,    2.65,    2.65,    2.65,
  2.46,    2.46,    2.46,    2.46,
  2.39,    2.39,    2.39,    2.39,
  2.21,    2.21,    2.21,    2.21,
  2.09,    2.09,    2.09,    2.09,
  1.9,     1.9,     1.9,     1.9,
  2.22,    2.22,    2.22,    2.22,
  2.34,    2.34,    2.34,    2.34,
  3.24,    3.24,    3.24,    3.24,
  3.45,    3.45,    3.45,    3.45,
  2.79,    2.79,    2.79,    2.79,
  2.8,     2.8,     2.8,     2.8,
  2.54,    2.54,    2.54,    2.54,
  2.24,    2.24,    2.24,    2.24,
  2.25,    2.25,    2.25,    2.25,
  1.91,    1.91,    1.91,    1.91,
  1.88,    1.88,    1.88,    1.88,
  1.87,    1.87,    1.87,    1.87,
  1.89,    1.89,    1.89,    1.89,
  1.59,    1.59,    1.59,    1.59,
  2.45,    2.45,    2.45,    2.45,
  2.14,    2.14,    2.14,    2.14,
  1.85,    1.85,    1.85,    1.85,
  1.77,    1.77,    1.77,    1.77,
  1.75,    1.75,    1.75,    1.75,
  1.29,    1.29,    1.29,    1.29,
  1.75,    1.75,    1.75,    1.75,
  1.26,    1.26,    1.26,    1.26,
  0.99,    0.99,    0.99,    0.99,
  0.69,    0.69,    0.69,    0.69,
  1,       1,       1,       1,
  0.84,    0.84,    0.84,    0.84,
  1.13,    1.13,    1.13,    1.13,
  0.77,    0.77,    0.77,    0.77,
  0.57,    0.57,    0.57,    0.57,
  0.64,    0.64,    0.64,    0.64,
  0.71,    0.71,    0.71,    0.71,
  1.48,    1.48,    1.48,    1.48,
  1.84,    1.84,    1.84,    1.84,
  1.55,    1.55,    1.55,    1.55,
  1.77,    1.77,    1.77,    1.77,
  1.62,    1.62,    1.62,    1.62,
  1.63,    1.63,    1.63,    1.63,
  1.55,    1.55,    1.55,    1.55,
  1.32,    1.32,    1.32,    1.32,
  1.52,    1.52,    1.52,    1.52,
  1.56,    1.56,    1.56,    1.56,
  1.16,    1.16,    1.16,    1.16,
  1.52,    1.52,    1.52,    1.52,
  1.65,    1.65,    1.65,    1.65,
  0.84,    0.84,    0.84,    0.84,
  0.96,    0.96,    0.96,    0.96,
  0.76,    0.76,    0.76,    0.76,
  0.18,    0.18,    0.18,    0.18,
  0.56,    0.56,    0.56,    0.56,
  0.61,    0.61,    0.61,    0.61,
  0.31,    0.31,    0.31,    0.31,
  0.31,    0.31,    0.31,    0.31,
  0.48,    0.48,    0.48,    0.48,
  0.62,    0.62,    0.62,    0.62,
  0.68,    0.68,    0.68,    0.68,
  0.54,    0.54,    0.54,    0.54,
  0.64,    0.64,    0.64,    0.64,
  0.79,    0.79,    0.79,    0.79,
  0.52,    0.52,    0.52,    0.52,
  0.94,    0.94,    0.94,    0.94,
  0.5,     0.5,     0.5,     0.5,
  1.22,    1.22,    1.22,    1.22,
  1.13,    1.13,    1.13,    1.13,
  0.64,    0.64,    0.64,    0.64,
  1.86,    1.86,    1.86,    1.86,
  1.85,    1.85,    1.85,    1.85,
  1.51,    1.51,    1.51,    1.51,
  1.48,    1.48,    1.48,    1.48,
  1.68,    1.68,    1.68,    1.68,
  1.83,    1.83,    1.83,    1.83,
  1.76,    1.76,    1.76,    1.76,
  1.16,    1.16,    1.16,    1.16,
  1.29,    1.29,    1.29,    1.29,
  1.67,    1.67,    1.67,    1.67,
  1.88,    1.88,    1.88,    1.88,
  1.69,    1.69,    1.69,    1.69,
  1.61,    1.61,    1.61,    1.61,
  1.53,    1.53,    1.53,    1.53,
  1.57,    1.57,    1.57,    1.57,
  1.5,     1.5,     1.5,     1.5,
  1.53,    1.53,    1.53,    1.53,
  1.36,    1.36,    1.36,    1.36,
  1.16,    1.16,    1.16,    1.16,
  1.23,    1.23,    1.23,    1.23,
  1.06,    1.06,    1.06,    1.06,
  0.92,    0.92,    0.92,    0.92,
  0.82,    0.82,    0.82,    0.82,
  1.02,    1.02,    1.02,    1.02,
  1.03,    1.03,    1.03,    1.03,
  0.79,    0.79,    0.79,    0.79,
  0.53,    0.53,    0.53,    0.53,
  0.87,    0.87,    0.87,    0.87,
  0.18,    0.18,    0.18,    0.18,
  0.1,     0.1,     0.1,     0.1,
  0.52,    0.52,    0.52,    0.52,
  0.42,    0.42,    0.42,    0.42,
  0.43,    0.43,    0.43,    0.43,
  0.64,    0.64,    0.64,    0.64,
  0.49,    0.49,    0.49,    0.49,
  0.76,    0.76,    0.76,    0.76,
  0.31,    0.31,    0.31,    0.31,
  0.66,    0.66,    0.66,    0.66,
  0.93,    0.93,    0.93,    0.93,
  0.1,     0.1,     0.1,     0.1,
  0.47,    0.47,    0.47,    0.47,
  0.1,     0.1,     0.1,     0.1,
  0.4,     0.4,     0.4,     0.4,
  0.04,    0.04,    0.04,    0.04,
  0.27,    0.27,    0.27,    0.27,
  0.84,    0.84,    0.84,    0.84,
  0.33,    0.33,    0.33,    0.33,
  0.36,    0.36,    0.36,    0.36,
  0.55,    0.55,    0.55,    0.55,
  0.19,    0.19,    0.19,    0.19,
  0.14,    0.14,    0.14,    0.14,
  0.28,    0.28,    0.28,    0.28,
  0.37,    0.37,    0.37,    0.37,
  1.71,    1.71,    1.71,    1.71,
  3.69,    3.69,    3.69,    3.69,
  4.34,    4.34,    4.34,    4.34,
  3.93,    3.93,    3.93,    3.93,
  4.03,    4.03,    4.03,    4.03,
  3.95,    3.95,    3.95,    3.95,
  3.42,    3.42,    3.42,    3.42,
  3.76,    3.76,    3.76,    3.76,
  3.33,    3.33,    3.33,    3.33,
  2.95,    2.95,    2.95,    2.95,
  3.22,    3.22,    3.22,    3.22,
  3.41,    3.41,    3.41,    3.41,
  3.31,    3.31,    3.31,    3.31,
  3.04,    3.04,    3.04,    3.04,
  3.14,    3.14,    3.14,    3.14,
  2.91,    2.91,    2.91,    2.91,
  3.04,    3.04,    3.04,    3.04,
  3.58,    3.58,    3.58,    3.58,
  3.9,     3.9,     3.9,     3.9,
  4.02,    4.02,    4.02,    4.02,
  4.22,    4.22,    4.22,    4.22,
  4.8,     4.8,     4.8,     4.8,
  4.59,    4.59,    4.59,    4.59,
  4.48,    4.48,    4.48,    4.48,
  4.47,    4.47,    4.47,    4.47,
  4.38,    4.38,    4.38,    4.38,
  4.46,    4.46,    4.46,    4.46,
  4.27,    4.27,    4.27,    4.27,
  4.32,    4.32,    4.32,    4.32,
  4.47,    4.47,    4.47,    4.47,
  4.67,    4.67,    4.67,    4.67,
  4.53,    4.53,    4.53,    4.53,
  3.91,    3.91,    3.91,    3.91,
  4.59,    4.59,    4.59,    4.59,
  4.71,    4.71,    4.71,    4.71,
  4.14,    4.14,    4.14,    4.14,
  4.16,    4.16,    4.16,    4.16,
  4.23,    4.23,    4.23,    4.23,
  3.8,     3.8,     3.8,     3.8,
  4.07,    4.07,    4.07,    4.07,
  4.26,    4.26,    4.26,    4.26,
  4.15,    4.15,    4.15,    4.15,
  4.17,    4.17,    4.17,    4.17,
  3.81,    3.81,    3.81,    3.81,
  3.63,    3.63,    3.63,    3.63,
  3.78,    3.78,    3.78,    3.78,
  3.86,    3.86,    3.86,    3.86,
  4.23,    4.23,    4.23,    4.23,
  4.6,     4.6,     4.6,     4.6,
  3.76,    3.76,    3.76,    3.76,
  4.15,    4.15,    4.15,    4.15,
  3.72,    3.72,    3.72,    3.72,
  4.05,    4.05,    4.05,    4.05,
  4,       4,       4,       4,
  4.44,    4.44,    4.44,    4.44,
  4.38,    4.38,    4.38,    4.38,
  4.13,    4.13,    4.13,    4.13,
  3.55,    3.55,    3.55,    3.55,
  3.01,    3.01,    3.01,    3.01,
  3.15,    3.15,    3.15,    3.15,
  3.48,    3.48,    3.48,    3.48,
  4.09,    4.09,    4.09,    4.09,
  3.82,    3.82,    3.82,    3.82,
  3.21,    3.21,    3.21,    3.21,
  3.31,    3.31,    3.31,    3.31,
  3.39,    3.39,    3.39,    3.39,
  3.34,    3.34,    3.34,    3.34,
  2.51,    2.51,    2.51,    2.51,
  2.83,    2.83,    2.83,    2.83,
  3.16,    3.16,    3.16,    3.16,
  2.93,    2.93,    2.93,    2.93,
  3.22,    3.22,    3.22,    3.22,
  3.16,    3.16,    3.16,    3.16,
  2.83,    2.83,    2.83,    2.83,
  2.72,    2.72,    2.72,    2.72,
  2.8,     2.8,     2.8,     2.8,
  3,       3,       3,       3,
  2.36,    2.36,    2.36,    2.36,
  2.31,    2.31,    2.31,    2.31,
  2.4,     2.4,     2.4,     2.4,
  2.4,     2.4,     2.4,     2.4,
  2.45,    2.45,    2.45,    2.45,
  2.16,    2.16,    2.16,    2.16,
  2.57,    2.57,    2.57,    2.57,
  2.96,    2.96,    2.96,    2.96,
  2.66,    2.66,    2.66,    2.66,
  2.75,    2.75,    2.75,    2.75,
  2.98,    2.98,    2.98,    2.98,
  2.71,    2.71,    2.71,    2.71,
  2.78,    2.78,    2.78,    2.78,
  2.73,    2.73,    2.73,    2.73,
  2.64,    2.64,    2.64,    2.64,
  2.61,    2.61,    2.61,    2.61,
  2.9,     2.9,     2.9,     2.9,
  2.77,    2.77,    2.77,    2.77,
  2.77,    2.77,    2.77,    2.77,
  3.36,    3.36,    3.36,    3.36,
  3.47,    3.47,    3.47,    3.47,
  2.76,    2.76,    2.76,    2.76,
  3.04,    3.04,    3.04,    3.04,
  3.31,    3.31,    3.31,    3.31,
  3.58,    3.58,    3.58,    3.58,
  3.1,     3.1,     3.1,     3.1,
  2.85,    2.85,    2.85,    2.85,
  2.58,    2.58,    2.58,    2.58,
  2.13,    2.13,    2.13,    2.13,
  2.6,     2.6,     2.6,     2.6,
  2.61,    2.61,    2.61,    2.61,
  2.71,    2.71,    2.71,    2.71,
  2.86,    2.86,    2.86,    2.86,
  2.63,    2.63,    2.63,    2.63,
  2.96,    2.96,    2.96,    2.96,
  2.9,     2.9,     2.9,     2.9,
  2.5,     2.5,     2.5,     2.5,
  2.62,    2.62,    2.62,    2.62,
  3.16,    3.16,    3.16,    3.16,
  3.42,    3.42,    3.42,    3.42,
  2.95,    2.95,    2.95,    2.95,
  3.04,    3.04,    3.04,    3.04,
  2.76,    2.76,    2.76,    2.76,
  2.77,    2.77,    2.77,    2.77,
  2.79,    2.79,    2.79,    2.79,
  3.03,    3.03,    3.03,    3.03,
  2.99,    2.99,    2.99,    2.99,
  3.1,     3.1,     3.1,     3.1,
  2.88,    2.88,    2.88,    2.88,
  2.54,    2.54,    2.54,    2.54,
  2.74,    2.74,    2.74,    2.74,
  3.14,    3.14,    3.14,    3.14,
  3.06,    3.06,    3.06,    3.06,
  2.98,    2.98,    2.98,    2.98,
  2.65,    2.65,    2.65,    2.65,
  2.54,    2.54,    2.54,    2.54,
  2.43,    2.43,    2.43,    2.43,
  2.33,    2.33,    2.33,    2.33,
  2.27,    2.27,    2.27,    2.27,
  2.46,    2.46,    2.46,    2.46,
  2.51,    2.51,    2.51,    2.51,
  2.39,    2.39,    2.39,    2.39,
  2.53,    2.53,    2.53,    2.53,
  2.65,    2.65,    2.65,    2.65,
  2.28,    2.28,    2.28,    2.28,
  2.87,    2.87,    2.87,    2.87,
  2.85,    2.85,    2.85,    2.85,
  3.12,    3.12,    3.12,    3.12,
  3.34,    3.34,    3.34,    3.34,
  3.12,    3.12,    3.12,    3.12,
  2.67,    2.67,    2.67,    2.67,
  2.88,    2.88,    2.88,    2.88,
  3.12,    3.12,    3.12,    3.12,
  3.03,    3.03,    3.03,    3.03,
  2.73,    2.73,    2.73,    2.73,
  2.9,     2.9,     2.9,     2.9,
  2.31,    2.31,    2.31,    2.31,
  2.16,    2.16,    2.16,    2.16,
  1.73,    1.73,    1.73,    1.73,
  1.98,    1.98,    1.98,    1.98,
  2.02,    2.02,    2.02,    2.02,
  2.06,    2.06,    2.06,    2.06,
  2,       2,       2,       2,
  1.97,    1.97,    1.97,    1.97,
  2.16,    2.16,    2.16,    2.16,
  2.17,    2.17,    2.17,    2.17,
  1.85,    1.85,    1.85,    1.85,
  1.69,    1.69,    1.69,    1.69,
  1.48,    1.48,    1.48,    1.48,
  2.51,    2.51,    2.51,    2.51,
  2.37,    2.37,    2.37,    2.37,
  2.38,    2.38,    2.38,    2.38,
  2.75,    2.75,    2.75,    2.75,
  2.83,    2.83,    2.83,    2.83,
  2.62,    2.62,    2.62,    2.62,
  3.32,    3.32,    3.32,    3.32,
  4.34,    4.34,    4.34,    4.34,
  3.36,    3.36,    3.36,    3.36,
  4.04,    4.04,    4.04,    4.04,
  4.29,    4.29,    4.29,    4.29,
  3.96,    3.96,    3.96,    3.96,
  3.45,    3.45,    3.45,    3.45,
  3.78,    3.78,    3.78,    3.78,
  3.47,    3.47,    3.47,    3.47,
  4,       4,       4,       4,
  5.76,    5.76,    5.76,    5.76,
  7.67,    7.67,    7.67,    7.67,
  6.78,    6.78,    6.78,    6.78,
  6.79,    6.79,    6.79,    6.79,
  5.59,    5.59,    5.59,    5.59,
  5.26,    5.26,    5.26,    5.26,
  4.98,    4.98,    4.98,    4.98,
  4.87,    4.87,    4.87,    4.87,
  5.02,    5.02,    5.02,    5.02,
  5.8,     5.8,     5.8,     5.8,
  5.69,    5.69,    5.69,    5.69,
  5.61,    5.61,    5.61,    5.61,
  5.48,    5.48,    5.48,    5.48,
  5.82,    5.82,    5.82,    5.82,
  5.6,     5.6,     5.6,     5.6,
  4.82,    4.82,    4.82,    4.82,
  4.72,    4.72,    4.72,    4.72,
  4.34,    4.34,    4.34,    4.34,
  4.27,    4.27,    4.27,    4.27,
  4.19,    4.19,    4.19,    4.19,
  4.31,    4.31,    4.31,    4.31,
  3.79,    3.79,    3.79,    3.79,
  3.86,    3.86,    3.86,    3.86,
  3.82,    3.82,    3.82,    3.82,
  3.99,    3.99,    3.99,    3.99,
  3.81,    3.81,    3.81,    3.81,
  3.43,    3.43,    3.43,    3.43,
  3.7,     3.7,     3.7,     3.7,
  3.48,    3.48,    3.48,    3.48,
  3.29,    3.29,    3.29,    3.29,
  3.39,    3.39,    3.39,    3.39,
  3.36,    3.36,    3.36,    3.36,
  3.06,    3.06,    3.06,    3.06,
  2.77,    2.77,    2.77,    2.77,
  2.63,    2.63,    2.63,    2.63,
  2.6,     2.6,     2.6,     2.6,
  2.7,     2.7,     2.7,     2.7,
  2.95,    2.95,    2.95,    2.95,
  2.9,     2.9,     2.9,     2.9,
  3.06,    3.06,    3.06,    3.06,
  2.8,     2.8,     2.8,     2.8,
  3.02,    3.02,    3.02,    3.02,
  2.9,     2.9,     2.9,     2.9,
  3,       3,       3,       3,
  3.44,    3.44,    3.44,    3.44,
  3.73,    3.73,    3.73,    3.73,
  3.98,    3.98,    3.98,    3.98,
  3.99,    3.99,    3.99,    3.99,
  3.87,    3.87,    3.87,    3.87,
  3.57,    3.57,    3.57,    3.57,
  3.42,    3.42,    3.42,    3.42,
  3.6,     3.6,     3.6,     3.6,
  3.44,    3.44,    3.44,    3.44,
  3.55,    3.55,    3.55,    3.55,
  4.1,     4.1,     4.1,     4.1,
  3.96,    3.96,    3.96,    3.96,
  4.1,     4.1,     4.1,     4.1,
  4.21,    4.21,    4.21,    4.21,
  4.28,    4.28,    4.28,    4.28,
  4.36,    4.36,    4.36,    4.36,
  4.26,    4.26,    4.26,    4.26,
  5.1,     5.1,     5.1,     5.1,
  4.9,     4.9,     4.9,     4.9,
  4.61,    4.61,    4.61,    4.61,
  4,       4,       4,       4,
  4.41,    4.41,    4.41,    4.41,
  4.49,    4.49,    4.49,    4.49,
  4.42,    4.42,    4.42,    4.42,
  3.75,    3.75,    3.75,    3.75,
  3.88,    3.88,    3.88,    3.88,
  3.7,     3.7,     3.7,     3.7,
  3.42,    3.42,    3.42,    3.42,
  3.16,    3.16,    3.16,    3.16,
  3.95,    3.95,    3.95,    3.95,
  3.84,    3.84,    3.84,    3.84,
  3.75,    3.75,    3.75,    3.75,
  3.6,     3.6,     3.6,     3.6,
  3.75,    3.75,    3.75,    3.75,
  4.17,    4.17,    4.17,    4.17,
  3.8,     3.8,     3.8,     3.8,
  3.69,    3.69,    3.69,    3.69,
  4.41,    4.41,    4.41,    4.41,
  4.84,    4.84,    4.84,    4.84,
  4.46,    4.46,    4.46,    4.46,
  4.53,    4.53,    4.53,    4.53,
  5.01,    5.01,    5.01,    5.01,
  4.46,    4.46,    4.46,    4.46,
  4.17,    4.17,    4.17,    4.17,
  3.82,    3.82,    3.82,    3.82,
  4.45,    4.45,    4.45,    4.45,
  4.28,    4.28,    4.28,    4.28,
  4.07,    4.07,    4.07,    4.07,
  3.86,    3.86,    3.86,    3.86,
  3.46,    3.46,    3.46,    3.46,
  3.38,    3.38,    3.38,    3.38,
  3.51,    3.51,    3.51,    3.51,
  3.39,    3.39,    3.39,    3.39,
  3.91,    3.91,    3.91,    3.91,
  3.24,    3.24,    3.24,    3.24,
  2.29,    2.29,    2.29,    2.29,
  2.53,    2.53,    2.53,    2.53,
  2.8,     2.8,     2.8,     2.8,
  3.04,    3.04,    3.04,    3.04,
  3.3,     3.3,     3.3,     3.3,
  3.89,    3.89,    3.89,    3.89,
  4.4,     4.4,     4.4,     4.4,
  4.5,     4.5,     4.5,     4.5,
  4.14,    4.14,    4.14,    4.14,
  4.66,    4.66,    4.66,    4.66,
  4.24,    4.24,    4.24,    4.24,
  4.59,    4.59,    4.59,    4.59,
  4.17,    4.17,    4.17,    4.17,
  4.59,    4.59,    4.59,    4.59,
  4.32,    4.32,    4.32,    4.32,
  3.82,    3.82,    3.82,    3.82,
  3.29,    3.29,    3.29,    3.29,
  3.06,    3.06,    3.06,    3.06,
  3.32,    3.32,    3.32,    3.32,
  3.4,     3.4,     3.4,     3.4,
  3.3,     3.3,     3.3,     3.3,
  3.77,    3.77,    3.77,    3.77,
  3.85,    3.85,    3.85,    3.85,
  3.73,    3.73,    3.73,    3.73,
  3.73,    3.73,    3.73,    3.73,
  3.8,     3.8,     3.8,     3.8,
  3.82,    3.82,    3.82,    3.82,
  3.44,    3.44,    3.44,    3.44,
  2.86,    2.86,    2.86,    2.86,
  2.78,    2.78,    2.78,    2.78,
  2.91,    2.91,    2.91,    2.91,
  2.8,     2.8,     2.8,     2.8,
  2.56,    2.56,    2.56,    2.56,
  3.45,    3.45,    3.45,    3.45,
  3.45,    3.45,    3.45,    3.45,
  2.97,    2.97,    2.97,    2.97,
  3.35,    3.35,    3.35,    3.35,
  2.85,    2.85,    2.85,    2.85,
  3.89,    3.89,    3.89,    3.89,
  4.09,    4.09,    4.09,    4.09,
  3.55,    3.55,    3.55,    3.55,
  3.29,    3.29,    3.29,    3.29,
  3.28,    3.28,    3.28,    3.28,
  3.46,    3.46,    3.46,    3.46,
  3.53,    3.53,    3.53,    3.53,
  3.37,    3.37,    3.37,    3.37,
  3.7,     3.7,     3.7,     3.7,
  3.31,    3.31,    3.31,    3.31,
  3.67,    3.67,    3.67,    3.67,
  3.8,     3.8,     3.8,     3.8,
  3.99,    3.99,    3.99,    3.99,
  3.33,    3.33,    3.33,    3.33,
  3.81,    3.81,    3.81,    3.81,
  4.31,    4.31,    4.31,    4.31,
  4.98,    4.98,    4.98,    4.98,
  4.38,    4.38,    4.38,    4.38,
  4.7,     4.7,     4.7,     4.7,
  4.85,    4.85,    4.85,    4.85,
  4.43,    4.43,    4.43,    4.43,
  4.02,    4.02,    4.02,    4.02,
  4.39,    4.39,    4.39,    4.39,
  3.62,    3.62,    3.62,    3.62,
  2.83,    2.83,    2.83,    2.83,
  2.83,    2.83,    2.83,    2.83,
  3.37,    3.37,    3.37,    3.37,
  3.7,     3.7,     3.7,     3.7,
  3.16,    3.16,    3.16,    3.16,
  3.49,    3.49,    3.49,    3.49,
  2.58,    2.58,    2.58,    2.58,
  3.01,    3.01,    3.01,    3.01,
  2.82,    2.82,    2.82,    2.82,
  2.69,    2.69,    2.69,    2.69,
  3.02,    3.02,    3.02,    3.02,
  3.27,    3.27,    3.27,    3.27,
  3.11,    3.11,    3.11,    3.11,
  3.27,    3.27,    3.27,    3.27,
  3.43,    3.43,    3.43,    3.43,
  3.66,    3.66,    3.66,    3.66,
  3.21,    3.21,    3.21,    3.21,
  3.05,    3.05,    3.05,    3.05,
  3.46,    3.46,    3.46,    3.46,
  3.22,    3.22,    3.22,    3.22,
  3.05,    3.05,    3.05,    3.05,
  3.75,    3.75,    3.75,    3.75,
  3.77,    3.77,    3.77,    3.77,
  3.63,    3.63,    3.63,    3.63,
  3.78,    3.78,    3.78,    3.78,
  4.02,    4.02,    4.02,    4.02,
  3.85,    3.85,    3.85,    3.85,
  4.11,    4.11,    4.11,    4.11,
  3.95,    3.95,    3.95,    3.95,
  3.47,    3.47,    3.47,    3.47,
  3.13,    3.13,    3.13,    3.13,
  3.27,    3.27,    3.27,    3.27,
  3.17,    3.17,    3.17,    3.17,
  3.07,    3.07,    3.07,    3.07,
  2.86,    2.86,    2.86,    2.86,
  2.9,     2.9,     2.9,     2.9,
  2.84,    2.84,    2.84,    2.84,
  3.44,    3.44,    3.44,    3.44,
  3.16,    3.16,    3.16,    3.16,
  3.06,    3.06,    3.06,    3.06,
  3.59,    3.59,    3.59,    3.59,
  3.18,    3.18,    3.18,    3.18,
  3.53,    3.53,    3.53,    3.53,
  3.79,    3.79,    3.79,    3.79,
  3.27,    3.27,    3.27,    3.27,
  2.95,    2.95,    2.95,    2.95,
  3.85,    3.85,    3.85,    3.85,
  3.4,     3.4,     3.4,     3.4,
  2.79,    2.79,    2.79,    2.79,
  2.55,    2.55,    2.55,    2.55,
  2.14,    2.14,    2.14,    2.14,
  1.91,    1.91,    1.91,    1.91,
  1.85,    1.85,    1.85,    1.85,
  1.74,    1.74,    1.74,    1.74,
  2.27,    2.27,    2.27,    2.27,
  2.27,    2.27,    2.27,    2.27,
  2.18,    2.18,    2.18,    2.18,
  1.92,    1.92,    1.92,    1.92,
  2.1,     2.1,     2.1,     2.1,
  2.03,    2.03,    2.03,    2.03,
  2.1,     2.1,     2.1,     2.1,
  2.19,    2.19,    2.19,    2.19,
  2.3,     2.3,     2.3,     2.3,
  2.48,    2.48,    2.48,    2.48,
  2.01,    2.01,    2.01,    2.01,
  1.67,    1.67,    1.67,    1.67,
  1.73,    1.73,    1.73,    1.73,
  2.11,    2.11,    2.11,    2.11,
  2.04,    2.04,    2.04,    2.04,
  2.24,    2.24,    2.24,    2.24,
  1.6,     1.6,     1.6,     1.6,
  1.23,    1.23,    1.23,    1.23,
  1.54,    1.54,    1.54,    1.54,
  1.75,    1.75,    1.75,    1.75,
  1.82,    1.82,    1.82,    1.82,
  1.38,    1.38,    1.38,    1.38,
  2.23,    2.23,    2.23,    2.23,
  2.14,    2.14,    2.14,    2.14,
  1.16,    1.16,    1.16,    1.16,
  0.8,     0.8,     0.8,     0.8,
  0.38,    0.38,    0.38,    0.38,
  1.35,    1.35,    1.35,    1.35,
  2.49,    2.49,    2.49,    2.49,
  1.88,    1.88,    1.88,    1.88,
  1.26,    1.26,    1.26,    1.26,
  1.45,    1.45,    1.45,    1.45,
  0.68,    0.68,    0.68,    0.68,
  0.35,    0.35,    0.35,    0.35,
  0.81,    0.81,    0.81,    0.81,
  0.72,    0.72,    0.72,    0.72,
  0.8,     0.8,     0.8,     0.8,
  0.94,    0.94,    0.94,    0.94,
  0.76,    0.76,    0.76,    0.76,
  1.26,    1.26,    1.26,    1.26,
  1.21,    1.21,    1.21,    1.21,
  0.81,    0.81,    0.81,    0.81,
  0.89,    0.89,    0.89,    0.89,
  0.92,    0.92,    0.92,    0.92,
  1.07,    1.07,    1.07,    1.07,
  1.53,    1.53,    1.53,    1.53,
  1.52,    1.52,    1.52,    1.52,
  1.17,    1.17,    1.17,    1.17,
  1.67,    1.67,    1.67,    1.67,
  2,       2,       2,       2,
  1.99,    1.99,    1.99,    1.99,
  1.76,    1.76,    1.76,    1.76,
  1.55,    1.55,    1.55,    1.55,
  1.15,    1.15,    1.15,    1.15,
  0.96,    0.96,    0.96,    0.96,
  1.51,    1.51,    1.51,    1.51,
  1.49,    1.49,    1.49,    1.49,
  1.82,    1.82,    1.82,    1.82,
  1.71,    1.71,    1.71,    1.71,
  1.59,    1.59,    1.59,    1.59,
  1.91,    1.91,    1.91,    1.91,
  1.98,    1.98,    1.98,    1.98,
  1.48,    1.48,    1.48,    1.48,
  1.62,    1.62,    1.62,    1.62,
  1.73,    1.73,    1.73,    1.73,
  1.41,    1.41,    1.41,    1.41,
  1.5,     1.5,     1.5,     1.5,
  1.29,    1.29,    1.29,    1.29,
  0.93,    0.93,    0.93,    0.93,
  1.38,    1.38,    1.38,    1.38,
  1.55,    1.55,    1.55,    1.55,
  1.37,    1.37,    1.37,    1.37,
  1.43,    1.43,    1.43,    1.43,
  1.26,    1.26,    1.26,    1.26,
  1.56,    1.56,    1.56,    1.56,
  1.52,    1.52,    1.52,    1.52,
  1.95,    1.95,    1.95,    1.95,
  2.04,    2.04,    2.04,    2.04,
  1.99,    1.99,    1.99,    1.99,
  2.22,    2.22,    2.22,    2.22,
  2.05,    2.05,    2.05,    2.05,
  2.27,    2.27,    2.27,    2.27,
  2.44,    2.44,    2.44,    2.44,
  2.32,    2.32,    2.32,    2.32,
  2.69,    2.69,    2.69,    2.69,
  2.8,     2.8,     2.8,     2.8,
  2.65,    2.65,    2.65,    2.65,
  2.12,    2.12,    2.12,    2.12,
  2.72,    2.72,    2.72,    2.72,
  2.43,    2.43,    2.43,    2.43,
  2.54,    2.54,    2.54,    2.54,
  2.28,    2.28,    2.28,    2.28,
  2.2,     2.2,     2.2,     2.2,
  2.19,    2.19,    2.19,    2.19,
  2.52,    2.52,    2.52,    2.52,
  2.87,    2.87,    2.87,    2.87,
  2.76,    2.76,    2.76,    2.76,
  2.51,    2.51,    2.51,    2.51,
  2.64,    2.64,    2.64,    2.64,
  2.12,    2.12,    2.12,    2.12,
  2.02,    2.02,    2.02,    2.02,
  1.98,    1.98,    1.98,    1.98,
  1.78,    1.78,    1.78,    1.78,
  2.2,     2.2,     2.2,     2.2,
  1.96,    1.96,    1.96,    1.96,
  1.54,    1.54,    1.54,    1.54,
  1.45,    1.45,    1.45,    1.45,
  1.7,     1.7,     1.7,     1.7,
  1.57,    1.57,    1.57,    1.57,
  1.5,     1.5,     1.5,     1.5,
  1.3,     1.3,     1.3,     1.3,
  1.92,    1.92,    1.92,    1.92,
  1.9,     1.9,     1.9,     1.9,
  1.44,    1.44,    1.44,    1.44,
  1.65,    1.65,    1.65,    1.65,
  1.72,    1.72,    1.72,    1.72,
  2.02,    2.02,    2.02,    2.02,
  1.85,    1.85,    1.85,    1.85,
  1.85,    1.85,    1.85,    1.85,
  2.06,    2.06,    2.06,    2.06,
  2.03,    2.03,    2.03,    2.03,
  2.23,    2.23,    2.23,    2.23,
  2.18,    2.18,    2.18,    2.18,
  2.23,    2.23,    2.23,    2.23,
  2.06,    2.06,    2.06,    2.06,
  2.22,    2.22,    2.22,    2.22,
  2.15,    2.15,    2.15,    2.15,
  2.15,    2.15,    2.15,    2.15,
  2.38,    2.38,    2.38,    2.38,
  2.46,    2.46,    2.46,    2.46,
  2.79,    2.79,    2.79,    2.79,
  2.54,    2.54,    2.54,    2.54,
  2.45,    2.45,    2.45,    2.45,
  2.96,    2.96,    2.96,    2.96,
  2.66,    2.66,    2.66,    2.66,
  2.24,    2.24,    2.24,    2.24,
  2.32,    2.32,    2.32,    2.32,
  2.71,    2.71,    2.71,    2.71,
  2.5,     2.5,     2.5,     2.5,
  1.99,    1.99,    1.99,    1.99,
  1.83,    1.83,    1.83,    1.83,
  1.91,    1.91,    1.91,    1.91,
  2.11,    2.11,    2.11,    2.11,
  2.15,    2.15,    2.15,    2.15,
  1.96,    1.96,    1.96,    1.96,
  2.33,    2.33,    2.33,    2.33,
  2.24,    2.24,    2.24,    2.24,
  2.38,    2.38,    2.38,    2.38,
  2.71,    2.71,    2.71,    2.71,
  2.07,    2.07,    2.07,    2.07,
  2.66,    2.66,    2.66,    2.66,
  2.84,    2.84,    2.84,    2.84,
  2.62,    2.62,    2.62,    2.62,
  3.22,    3.22,    3.22,    3.22,
  3.32,    3.32,    3.32,    3.32,
  3.69,    3.69,    3.69,    3.69,
  3.69,    3.69,    3.69,    3.69,
  3.48,    3.48,    3.48,    3.48,
  3.43,    3.43,    3.43,    3.43,
  3.83,    3.83,    3.83,    3.83,
  3.63,    3.63,    3.63,    3.63,
  3.63,    3.63,    3.63,    3.63,
  3.53,    3.53,    3.53,    3.53,
  3.4,     3.4,     3.4,     3.4,
  3.34,    3.34,    3.34,    3.34,
  2.94,    2.94,    2.94,    2.94,
  3.23,    3.23,    3.23,    3.23,
  3.29,    3.29,    3.29,    3.29,
  3.16,    3.16,    3.16,    3.16,
  2.66,    2.66,    2.66,    2.66,
  2.7,     2.7,     2.7,     2.7,
  2.87,    2.87,    2.87,    2.87,
  2.33,    2.33,    2.33,    2.33,
  2.36,    2.36,    2.36,    2.36,
  2.11,    2.11,    2.11,    2.11,
  2.29,    2.29,    2.29,    2.29,
  2.36,    2.36,    2.36,    2.36,
  2.02,    2.02,    2.02,    2.02,
  2.47,    2.47,    2.47,    2.47,
  2.5,     2.5,     2.5,     2.5,
  2.61,    2.61,    2.61,    2.61,
  2.12,    2.12,    2.12,    2.12,
  2.23,    2.23,    2.23,    2.23,
  2.03,    2.03,    2.03,    2.03,
  2.13,    2.13,    2.13,    2.13,
  2.41,    2.41,    2.41,    2.41,
  2.8,     2.8,     2.8,     2.8,
  2.47,    2.47,    2.47,    2.47,
  2.44,    2.44,    2.44,    2.44,
  1.69,    1.69,    1.69,    1.69,
  1.75,    1.75,    1.75,    1.75,
  1.92,    1.92,    1.92,    1.92,
  2.05,    2.05,    2.05,    2.05,
  1.82,    1.82,    1.82,    1.82,
  2.09,    2.09,    2.09,    2.09,
  1.57,    1.57,    1.57,    1.57,
  1.62,    1.62,    1.62,    1.62,
  1.88,    1.88,    1.88,    1.88,
  1.74,    1.74,    1.74,    1.74,
  1.99,    1.99,    1.99,    1.99,
  1.61,    1.61,    1.61,    1.61,
  1.36,    1.36,    1.36,    1.36,
  1.38,    1.38,    1.38,    1.38,
  1.78,    1.78,    1.78,    1.78,
  1.53,    1.53,    1.53,    1.53,
  0.85,    0.85,    0.85,    0.85,
  0.78,    0.78,    0.78,    0.78,
  1.06,    1.06,    1.06,    1.06,
  0.92,    0.92,    0.92,    0.92,
  1.22,    1.22,    1.22,    1.22,
  1.19,    1.19,    1.19,    1.19,
  1.29,    1.29,    1.29,    1.29,
  1.18,    1.18,    1.18,    1.18,
  1.19,    1.19,    1.19,    1.19,
  1.48,    1.48,    1.48,    1.48,
  1.9,     1.9,     1.9,     1.9,
  1.68,    1.68,    1.68,    1.68,
  1.4,     1.4,     1.4,     1.4,
  1.47,    1.47,    1.47,    1.47,
  1.34,    1.34,    1.34,    1.34,
  2.04,    2.04,    2.04,    2.04,
  1.92,    1.92,    1.92,    1.92,
  2.12,    2.12,    2.12,    2.12,
  2.71,    2.71,    2.71,    2.71,
  2.11,    2.11,    2.11,    2.11,
  2.54,    2.54,    2.54,    2.54,
  2.29,    2.29,    2.29,    2.29,
  2.37,    2.37,    2.37,    2.37,
  2.31,    2.31,    2.31,    2.31,
  2.45,    2.45,    2.45,    2.45,
  2.28,    2.28,    2.28,    2.28,
  2.57,    2.57,    2.57,    2.57,
  2.44,    2.44,    2.44,    2.44,
  2.57,    2.57,    2.57,    2.57,
  2.95,    2.95,    2.95,    2.95,
  2.8,     2.8,     2.8,     2.8,
  2.66,    2.66,    2.66,    2.66,
  2.71,    2.71,    2.71,    2.71,
  2.58,    2.58,    2.58,    2.58,
  2.94,    2.94,    2.94,    2.94,
  2.61,    2.61,    2.61,    2.61,
  2.5,     2.5,     2.5,     2.5,
  2.97,    2.97,    2.97,    2.97,
  3.65,    3.65,    3.65,    3.65,
  3.56,    3.56,    3.56,    3.56,
  3.24,    3.24,    3.24,    3.24,
  3.35,    3.35,    3.35,    3.35,
  2.87,    2.87,    2.87,    2.87,
  2.85,    2.85,    2.85,    2.85,
  3.59,    3.59,    3.59,    3.59,
  3.14,    3.14,    3.14,    3.14,
  2.69,    2.69,    2.69,    2.69,
  2.28,    2.28,    2.28,    2.28,
  2.58,    2.58,    2.58,    2.58,
  2.61,    2.61,    2.61,    2.61,
  2.36,    2.36,    2.36,    2.36,
  2.64,    2.64,    2.64,    2.64,
  3.43,    3.43,    3.43,    3.43,
  3.22,    3.22,    3.22,    3.22,
  2.72,    2.72,    2.72,    2.72,
  2.8,     2.8,     2.8,     2.8,
  2.88,    2.88,    2.88,    2.88,
  3.01,    3.01,    3.01,    3.01,
  2.63,    2.63,    2.63,    2.63,
  2.63,    2.63,    2.63,    2.63,
  2.55,    2.55,    2.55,    2.55,
  2.44,    2.44,    2.44,    2.44,
  2.92,    2.92,    2.92,    2.92,
  3.23,    3.23,    3.23,    3.23,
  2.76,    2.76,    2.76,    2.76,
  3.12,    3.12,    3.12,    3.12,
  3.02,    3.02,    3.02,    3.02,
  3.51,    3.51,    3.51,    3.51,
  3.43,    3.43,    3.43,    3.43,
  4.18,    4.18,    4.18,    4.18,
  3.77,    3.77,    3.77,    3.77,
  4.12,    4.12,    4.12,    4.12,
  3.92,    3.92,    3.92,    3.92,
  3.95,    3.95,    3.95,    3.95,
  3.28,    3.28,    3.28,    3.28,
  3.36,    3.36,    3.36,    3.36,
  3.41,    3.41,    3.41,    3.41,
  3.32,    3.32,    3.32,    3.32,
  3.3,     3.3,     3.3,     3.3,
  3.15,    3.15,    3.15,    3.15,
  3.77,    3.77,    3.77,    3.77,
  3.7,     3.7,     3.7,     3.7,
  4.09,    4.09,    4.09,    4.09,
  3.43,    3.43,    3.43,    3.43,
  2.91,    2.91,    2.91,    2.91,
  2.39,    2.39,    2.39,    2.39,
  2.5,     2.5,     2.5,     2.5,
  2.59,    2.59,    2.59,    2.59,
  2.87,    2.87,    2.87,    2.87,
  3.34,    3.34,    3.34,    3.34,
  3.09,    3.09,    3.09,    3.09,
  3.69,    3.69,    3.69,    3.69,
  3.96,    3.96,    3.96,    3.96,
  3.89,    3.89,    3.89,    3.89,
  4.09,    4.09,    4.09,    4.09,
  3.38,    3.38,    3.38,    3.38,
  3.08,    3.08,    3.08,    3.08,
  3.68,    3.68,    3.68,    3.68,
  3.23,    3.23,    3.23,    3.23,
  3.4,     3.4,     3.4,     3.4,
  3.49,    3.49,    3.49,    3.49,
  3.46,    3.46,    3.46,    3.46,
  3.24,    3.24,    3.24,    3.24,
  3.07,    3.07,    3.07,    3.07,
  3.7,     3.7,     3.7,     3.7,
  3.68,    3.68,    3.68,    3.68,
  3.37,    3.37,    3.37,    3.37,
  3.25,    3.25,    3.25,    3.25,
  3.18,    3.18,    3.18,    3.18,
  3.44,    3.44,    3.44,    3.44,
  3.2,     3.2,     3.2,     3.2,
  3.29,    3.29,    3.29,    3.29,
  3.28,    3.28,    3.28,    3.28,
  3.92,    3.92,    3.92,    3.92,
  3.97,    3.97,    3.97,    3.97,
  5.2,     5.2,     5.2,     5.2,
  4.96,    4.96,    4.96,    4.96,
  4.93,    4.93,    4.93,    4.93,
  5.37,    5.37,    5.37,    5.37,
  4.84,    4.84,    4.84,    4.84,
  4.66,    4.66,    4.66,    4.66,
  4.93,    4.93,    4.93,    4.93,
  4.23,    4.23,    4.23,    4.23,
  4.56,    4.56,    4.56,    4.56,
  4.34,    4.34,    4.34,    4.34,
  4,       4,       4,       4,
  4,       4,       4,       4,
  3.64,    3.64,    3.64,    3.64,
  3.37,    3.37,    3.37,    3.37,
  3.34,    3.34,    3.34,    3.34,
  3.59,    3.59,    3.59,    3.59,
  3.66,    3.66,    3.66,    3.66,
  3.78,    3.78,    3.78,    3.78,
  3.46,    3.46,    3.46,    3.46,
  3.07,    3.07,    3.07,    3.07,
  2.86,    2.86,    2.86,    2.86,
  2.84,    2.84,    2.84,    2.84,
  3.13,    3.13,    3.13,    3.13,
  3.15,    3.15,    3.15,    3.15,
  3.55,    3.55,    3.55,    3.55,
  3.41,    3.41,    3.41,    3.41,
  3.32,    3.32,    3.32,    3.32,
  3.42,    3.42,    3.42,    3.42,
  3.57,    3.57,    3.57,    3.57,
  3.73,    3.73,    3.73,    3.73,
  3.38,    3.38,    3.38,    3.38,
  3.58,    3.58,    3.58,    3.58,
  3.58,    3.58,    3.58,    3.58,
  3.59,    3.59,    3.59,    3.59,
  3.47,    3.47,    3.47,    3.47,
  3.96,    3.96,    3.96,    3.96,
  3.5,     3.5,     3.5,     3.5,
  3.14,    3.14,    3.14,    3.14,
  2.81,    2.81,    2.81,    2.81,
  3.26,    3.26,    3.26,    3.26,
  3.65,    3.65,    3.65,    3.65,
  3.73,    3.73,    3.73,    3.73,
  3.77,    3.77,    3.77,    3.77,
  4.02,    4.02,    4.02,    4.02,
  3.92,    3.92,    3.92,    3.92,
  3.98,    3.98,    3.98,    3.98,
  3.88,    3.88,    3.88,    3.88,
  4.63,    4.63,    4.63,    4.63,
  4.46,    4.46,    4.46,    4.46,
  4.72,    4.72,    4.72,    4.72,
  4.67,    4.67,    4.67,    4.67,
  3.44,    3.44,    3.44,    3.44,
  4.13,    4.13,    4.13,    4.13,
  4.65,    4.65,    4.65,    4.65,
  4.78,    4.78,    4.78,    4.78,
  4.1,     4.1,     4.1,     4.1,
  4.73,    4.73,    4.73,    4.73,
  4.64,    4.64,    4.64,    4.64,
  4.36,    4.36,    4.36,    4.36,
  4.03,    4.03,    4.03,    4.03,
  3.17,    3.17,    3.17,    3.17,
  3.38,    3.38,    3.38,    3.38,
  3.08,    3.08,    3.08,    3.08,
  3.34,    3.34,    3.34,    3.34,
  4.2,     4.2,     4.2,     4.2,
  4.32,    4.32,    4.32,    4.32,
  3.91,    3.91,    3.91,    3.91,
  3.78,    3.78,    3.78,    3.78,
  3.59,    3.59,    3.59,    3.59,
  3.91,    3.91,    3.91,    3.91,
  3.17,    3.17,    3.17,    3.17,
  3.61,    3.61,    3.61,    3.61,
  3.17,    3.17,    3.17,    3.17,
  3.63,    3.63,    3.63,    3.63,
  3.91,    3.91,    3.91,    3.91,
  3.71,    3.71,    3.71,    3.71,
  3.26,    3.26,    3.26,    3.26,
  4.35,    4.35,    4.35,    4.35,
  4.22,    4.22,    4.22,    4.22,
  4,       4,       4,       4,
  3.57,    3.57,    3.57,    3.57,
  3.63,    3.63,    3.63,    3.63,
  3.47,    3.47,    3.47,    3.47,
  3.3,     3.3,     3.3,     3.3,
  3.5,     3.5,     3.5,     3.5,
  3.46,    3.46,    3.46,    3.46,
  3.77,    3.77,    3.77,    3.77,
  3.31,    3.31,    3.31,    3.31,
  3.65,    3.65,    3.65,    3.65,
  3.72,    3.72,    3.72,    3.72,
  4.37,    4.37,    4.37,    4.37,
  3.61,    3.61,    3.61,    3.61,
  3.81,    3.81,    3.81,    3.81,
  2.94,    2.94,    2.94,    2.94,
  3.15,    3.15,    3.15,    3.15,
  3.84,    3.84,    3.84,    3.84,
  3.48,    3.48,    3.48,    3.48,
  2.93,    2.93,    2.93,    2.93,
  3.77,    3.77,    3.77,    3.77,
  3.28,    3.28,    3.28,    3.28,
  4.02,    4.02,    4.02,    4.02,
  3.45,    3.45,    3.45,    3.45,
  3.42,    3.42,    3.42,    3.42,
  3.19,    3.19,    3.19,    3.19,
  3.59,    3.59,    3.59,    3.59,
  3.75,    3.75,    3.75,    3.75,
  3.53,    3.53,    3.53,    3.53,
  3.62,    3.62,    3.62,    3.62,
  3.98,    3.98,    3.98,    3.98,
  3.44,    3.44,    3.44,    3.44,
  3.46,    3.46,    3.46,    3.46,
  3.91,    3.91,    3.91,    3.91,
  3.86,    3.86,    3.86,    3.86,
  4.07,    4.07,    4.07,    4.07,
  4.01,    4.01,    4.01,    4.01,
  3.73,    3.73,    3.73,    3.73,
  3.61,    3.61,    3.61,    3.61,
  3.29,    3.29,    3.29,    3.29,
  3.42,    3.42,    3.42,    3.42,
  3.24,    3.24,    3.24,    3.24,
  3.58,    3.58,    3.58,    3.58,
  3.04,    3.04,    3.04,    3.04,
  3,       3,       3,       3,
  2.86,    2.86,    2.86,    2.86,
  2.67,    2.67,    2.67,    2.67,
  2.64,    2.64,    2.64,    2.64,
  2.43,    2.43,    2.43,    2.43,
  2.81,    2.81,    2.81,    2.81,
  2.98,    2.98,    2.98,    2.98,
  2.5,     2.5,     2.5,     2.5,
  3.08,    3.08,    3.08,    3.08,
  3.27,    3.27,    3.27,    3.27,
  2.51,    2.51,    2.51,    2.51,
  2.11,    2.11,    2.11,    2.11,
  2.13,    2.13,    2.13,    2.13,
  2.16,    2.16,    2.16,    2.16,
  2.24,    2.24,    2.24,    2.24,
  1.97,    1.97,    1.97,    1.97,
  1.87,    1.87,    1.87,    1.87,
  2.21,    2.21,    2.21,    2.21,
  2,       2,       2,       2,
  2.05,    2.05,    2.05,    2.05,
  1.96,    1.96,    1.96,    1.96,
  2.02,    2.02,    2.02,    2.02,
  2.16,    2.16,    2.16,    2.16,
  2.47,    2.47,    2.47,    2.47,
  2.16,    2.16,    2.16,    2.16,
  2.21,    2.21,    2.21,    2.21,
  2.12,    2.12,    2.12,    2.12,
  2.19,    2.19,    2.19,    2.19,
  2.69,    2.69,    2.69,    2.69,
  1.68,    1.68,    1.68,    1.68,
  1.56,    1.56,    1.56,    1.56,
  1.1,     1.1,     1.1,     1.1,
  2.91,    2.91,    2.91,    2.91,
  2.978,   2.978,   2.978,   2.978,
  2.89,    2.89,    2.89,    2.89,
  2.988,   2.988,   2.988,   2.988,
  2.92,    2.92,    2.92,    2.92,
  3.02,    3.02,    3.02,    3.02,
  3.198,   3.198,   3.198,   3.198,
  3.18,    3.18,    3.18,    3.18,
  3.221,   3.221,   3.221,   3.221,
  3.145,   3.145,   3.145,   3.145,
  3.204,   3.204,   3.204,   3.204,
  3.208,   3.208,   3.208,   3.208,
  3.074,   3.074,   3.074,   3.074,
  3.036,   3.036,   3.036,   3.036,
  2.927,   2.927,   2.927,   2.927,
  2.81,    2.81,    2.81,    2.81,
  2.818,   2.818,   2.818,   2.818,
  2.921,   2.921,   2.921,   2.921,
  2.986,   2.986,   2.986,   2.986,
  3.054,   3.054,   3.054,   3.054,
  2.815,   2.815,   2.815,   2.815,
  2.823,   2.823,   2.823,   2.823,
  2.938,   2.938,   2.938,   2.938,
  2.879,   2.879,   2.879,   2.879,
  2.871,   2.871,   2.871,   2.871,
  2.991,   2.991,   2.991,   2.991,
  2.901,   2.901,   2.901,   2.901,
  2.82,    2.82,    2.82,    2.82,
  2.827,   2.827,   2.827,   2.827,
  2.776,   2.776,   2.776,   2.776,
  2.796,   2.796,   2.796,   2.796,
  2.741,   2.741,   2.741,   2.741,
  2.851,   2.851,   2.851,   2.851,
  2.806,   2.806,   2.806,   2.806,
  2.779,   2.779,   2.779,   2.779,
  2.738,   2.738,   2.738,   2.738,
  2.87,    2.87,    2.87,    2.87,
  3.034,   3.034,   3.034,   3.034,
  2.918,   2.918,   2.918,   2.918,
  2.93,    2.93,    2.93,    2.93,
  2.983,   2.983,   2.983,   2.983,
  2.696,   2.696,   2.696,   2.696,
  2.785,   2.785,   2.785,   2.785,
  2.815,   2.815,   2.815,   2.815,
  2.924,   2.924,   2.924,   2.924,
  2.685,   2.685,   2.685,   2.685,
  2.669,   2.669,   2.669,   2.669,
  2.763,   2.763,   2.763,   2.763,
  2.91,    2.91,    2.91,    2.91,
  2.978,   2.978,   2.978,   2.978,
  2.89,    2.89,    2.89,    2.89,
  2.988,   2.988,   2.988,   2.988,
  2.92,    2.92,    2.92,    2.92,
  3.02,    3.02,    3.02,    3.02,
  3.198,   3.198,   3.198,   3.198,
  3.18,    3.18,    3.18,    3.18,
  3.221,   3.221,   3.221,   3.221,
  3.145,   3.145,   3.145,   3.145,
  3.204,   3.204,   3.204,   3.204,
  3.208,   3.208,   3.208,   3.208,
  3.074,   3.074,   3.074,   3.074,
  3.036,   3.036,   3.036,   3.036,
  2.927,   2.927,   2.927,   2.927,
  2.81,    2.81,    2.81,    2.81,
  2.818,   2.818,   2.818,   2.818,
  2.921,   2.921,   2.921,   2.921,
  2.986,   2.986,   2.986,   2.986,
  3.054,   3.054,   3.054,   3.054,
  2.815,   2.815,   2.815,   2.815,
  2.823,   2.823,   2.823,   2.823,
  2.938,   2.938,   2.938,   2.938,
  2.879,   2.879,   2.879,   2.879,
  2.871,   2.871,   2.871,   2.871,
  2.991,   2.991,   2.991,   2.991,
  2.901,   2.901,   2.901,   2.901,
  2.82,    2.82,    2.82,    2.82,
  2.827,   2.827,   2.827,   2.827,
  2.776,   2.776,   2.776,   2.776,
  2.796,   2.796,   2.796,   2.796,
  2.741,   2.741,   2.741,   2.741,
  2.851,   2.851,   2.851,   2.851,
  2.806,   2.806,   2.806,   2.806,
  2.779,   2.779,   2.779,   2.779,
  2.738,   2.738,   2.738,   2.738,
  2.87,    2.87,    2.87,    2.87,
  3.034,   3.034,   3.034,   3.034,
  2.918,   2.918,   2.918,   2.918,
  2.93,    2.93,    2.93,    2.93,
  2.983,   2.983,   2.983,   2.983,
  2.696,   2.696,   2.696,   2.696,
  2.785,   2.785,   2.785,   2.785,
  2.815,   2.815,   2.815,   2.815,
  2.924,   2.924,   2.924,   2.924,
  2.685,   2.685,   2.685,   2.685,
  2.669,   2.669,   2.669,   2.669,
  2.763,   2.763,   2.763,   2.763,
  2.91,    2.91,    2.91,    2.91,
  2.978,   2.978,   2.978,   2.978,
  2.89,    2.89,    2.89,    2.89,
  2.988,   2.988,   2.988,   2.988,
  2.92,    2.92,    2.92,    2.92,
  3.02,    3.02,    3.02,    3.02,
  3.198,   3.198,   3.198,   3.198,
  3.18,    3.18,    3.18,    3.18,
  3.221,   3.221,   3.221,   3.221,
  3.145,   3.145,   3.145,   3.145,
  3.204,   3.204,   3.204,   3.204,
  3.208,   3.208,   3.208,   3.208,
  3.074,   3.074,   3.074,   3.074,
  3.036,   3.036,   3.036,   3.036,
  2.927,   2.927,   2.927,   2.927,
  2.81,    2.81,    2.81,    2.81,
  2.818,   2.818,   2.818,   2.818,
  2.921,   2.921,   2.921,   2.921,
  2.986,   2.986,   2.986,   2.986,
  3.054,   3.054,   3.054,   3.054,
  2.815,   2.815,   2.815,   2.815,
  2.823,   2.823,   2.823,   2.823,
  2.938,   2.938,   2.938,   2.938,
  2.879,   2.879,   2.879,   2.879,
  2.871,   2.871,   2.871,   2.871,
  2.991,   2.991,   2.991,   2.991,
  2.901,   2.901,   2.901,   2.901,
  2.82,    2.82,    2.82,    2.82,
  2.827,   2.827,   2.827,   2.827,
  2.776,   2.776,   2.776,   2.776,
  2.796,   2.796,   2.796,   2.796,
  2.741,   2.741,   2.741,   2.741,
  2.851,   2.851,   2.851,   2.851,
  2.806,   2.806,   2.806,   2.806,
  2.779,   2.779,   2.779,   2.779,
  2.738,   2.738,   2.738,   2.738,
  2.87,    2.87,    2.87,    2.87,
  3.034,   3.034,   3.034,   3.034,
  2.918,   2.918,   2.918,   2.918,
  2.93,    2.93,    2.93,    2.93,
  2.983,   2.983,   2.983,   2.983,
  2.696,   2.696,   2.696,   2.696,
  2.785,   2.785,   2.785,   2.785,
  2.815,   2.815,   2.815,   2.815,
  2.924,   2.924,   2.924,   2.924,
  2.685,   2.685,   2.685,   2.685,
  2.669,   2.669,   2.669,   2.669,
  2.763,   2.763,   2.763,   2.763,
  3.29,    3.29,    3.29,    3.29,
  2.88,    2.88,    2.88,    2.88,
  2.57,    2.57,    2.57,    2.57,
  2.99,    2.99,    2.99,    2.99,
  2.96,    2.96,    2.96,    2.96,
  3.31,    3.31,    3.31,    3.31,
  3.16,    3.16,    3.16,    3.16,
  3.04,    3.04,    3.04,    3.04,
  3.2,     3.2,     3.2,     3.2,
  3.32,    3.32,    3.32,    3.32,
  3.68,    3.68,    3.68,    3.68,
  3.28,    3.28,    3.28,    3.28,
  3.38,    3.38,    3.38,    3.38,
  3.52,    3.52,    3.52,    3.52,
  3.61,    3.61,    3.61,    3.61,
  3.91,    3.91,    3.91,    3.91,
  3.69,    3.69,    3.69,    3.69,
  3.89,    3.89,    3.89,    3.89,
  3.72,    3.72,    3.72,    3.72,
  3.67,    3.67,    3.67,    3.67,
  3.43,    3.43,    3.43,    3.43,
  3.55,    3.55,    3.55,    3.55,
  3.5,     3.5,     3.5,     3.5,
  3.28,    3.28,    3.28,    3.28,
  3.26,    3.26,    3.26,    3.26,
  3.74,    3.74,    3.74,    3.74,
  3.76,    3.76,    3.76,    3.76,
  3.84,    3.84,    3.84,    3.84,
  3.72,    3.72,    3.72,    3.72,
  2.98,    2.98,    2.98,    2.98,
  3.24,    3.24,    3.24,    3.24,
  3.03,    3.03,    3.03,    3.03,
  3.17,    3.17,    3.17,    3.17,
  3.32,    3.32,    3.32,    3.32,
  3.16,    3.16,    3.16,    3.16,
  3.09,    3.09,    3.09,    3.09,
  3.04,    3.04,    3.04,    3.04,
  3.22,    3.22,    3.22,    3.22,
  3.08,    3.08,    3.08,    3.08,
  3.17,    3.17,    3.17,    3.17,
  3.4,     3.4,     3.4,     3.4,
  3.06,    3.06,    3.06,    3.06,
  3.1,     3.1,     3.1,     3.1,
  2.79,    2.79,    2.79,    2.79,
  2.62,    2.62,    2.62,    2.62,
  3.27,    3.27,    3.27,    3.27,
  3.13,    3.13,    3.13,    3.13,
  2.89,    2.89,    2.89,    2.89,
  2.78,    2.78,    2.78,    2.78,
  2.95,    2.95,    2.95,    2.95,
  3.01,    3.01,    3.01,    3.01,
  2.95,    2.95,    2.95,    2.95,
  2.84,    2.84,    2.84,    2.84,
  2.96,    2.96,    2.96,    2.96,
  2.93,    2.93,    2.93,    2.93,
  3.35,    3.35,    3.35,    3.35,
  3.24,    3.24,    3.24,    3.24,
  3.2,     3.2,     3.2,     3.2,
  2.96,    2.96,    2.96,    2.96,
  2.85,    2.85,    2.85,    2.85,
  2.83,    2.83,    2.83,    2.83,
  2.82,    2.82,    2.82,    2.82,
  2.43,    2.43,    2.43,    2.43,
  2.11,    2.11,    2.11,    2.11,
  2.62,    2.62,    2.62,    2.62,
  2.71,    2.71,    2.71,    2.71,
  3.08,    3.08,    3.08,    3.08,
  3.63,    3.63,    3.63,    3.63,
  3.06,    3.06,    3.06,    3.06,
  3.29,    3.29,    3.29,    3.29,
  3.24,    3.24,    3.24,    3.24,
  2.77,    2.77,    2.77,    2.77,
  2.95,    2.95,    2.95,    2.95,
  3.05,    3.05,    3.05,    3.05,
  2.69,    2.69,    2.69,    2.69,
  3.18,    3.18,    3.18,    3.18,
  3.55,    3.55,    3.55,    3.55,
  3.73,    3.73,    3.73,    3.73,
  3.55,    3.55,    3.55,    3.55,
  4.19,    4.19,    4.19,    4.19,
  3.73,    3.73,    3.73,    3.73,
  3.27,    3.27,    3.27,    3.27,
  3.76,    3.76,    3.76,    3.76,
  3.96,    3.96,    3.96,    3.96,
  4.1,     4.1,     4.1,     4.1,
  4.12,    4.12,    4.12,    4.12,
  3.89,    3.89,    3.89,    3.89,
  4.05,    4.05,    4.05,    4.05,
  3.44,    3.44,    3.44,    3.44,
  3.66,    3.66,    3.66,    3.66,
  3.91,    3.91,    3.91,    3.91,
  3.65,    3.65,    3.65,    3.65,
  3.35,    3.35,    3.35,    3.35,
  3.85,    3.85,    3.85,    3.85,
  3.82,    3.82,    3.82,    3.82,
  4.33,    4.33,    4.33,    4.33,
  4.33,    4.33,    4.33,    4.33,
  5.14,    5.14,    5.14,    5.14,
  4.83,    4.83,    4.83,    4.83,
  4.73,    4.73,    4.73,    4.73,
  4.3,     4.3,     4.3,     4.3,
  4.3,     4.3,     4.3,     4.3,
  4.64,    4.64,    4.64,    4.64,
  4.27,    4.27,    4.27,    4.27,
  4.24,    4.24,    4.24,    4.24,
  4.12,    4.12,    4.12,    4.12,
  3.32,    3.32,    3.32,    3.32,
  4.24,    4.24,    4.24,    4.24,
  4.17,    4.17,    4.17,    4.17,
  3.69,    3.69,    3.69,    3.69,
  3.9,     3.9,     3.9,     3.9,
  3.85,    3.85,    3.85,    3.85,
  4.18,    4.18,    4.18,    4.18,
  4.27,    4.27,    4.27,    4.27,
  3.99,    3.99,    3.99,    3.99,
  3.76,    3.76,    3.76,    3.76,
  2.83,    2.83,    2.83,    2.83,
  3.08,    3.08,    3.08,    3.08,
  3.33,    3.33,    3.33,    3.33,
  3.67,    3.67,    3.67,    3.67,
  3.32,    3.32,    3.32,    3.32,
  3.14,    3.14,    3.14,    3.14,
  3.16,    3.16,    3.16,    3.16,
  3.17,    3.17,    3.17,    3.17,
  3.35,    3.35,    3.35,    3.35,
  2.81,    2.81,    2.81,    2.81,
  3.18,    3.18,    3.18,    3.18,
  3.38,    3.38,    3.38,    3.38,
  3.61,    3.61,    3.61,    3.61,
  3.87,    3.87,    3.87,    3.87,
  2.98,    2.98,    2.98,    2.98,
  2.18,    2.18,    2.18,    2.18,
  3.25,    3.25,    3.25,    3.25,
  3.31,    3.31,    3.31,    3.31,
  3.23,    3.23,    3.23,    3.23,
  3.22,    3.22,    3.22,    3.22,
  2.78,    2.78,    2.78,    2.78,
  3.23,    3.23,    3.23,    3.23,
  2.57,    2.57,    2.57,    2.57,
  2.91,    2.91,    2.91,    2.91,
  3.07,    3.07,    3.07,    3.07,
  2.31,    2.31,    2.31,    2.31,
  2.53,    2.53,    2.53,    2.53,
  2.78,    2.78,    2.78,    2.78,
  2.87,    2.87,    2.87,    2.87,
  3.2,     3.2,     3.2,     3.2,
  3.61,    3.61,    3.61,    3.61,
  3.49,    3.49,    3.49,    3.49,
  3.33,    3.33,    3.33,    3.33,
  3.19,    3.19,    3.19,    3.19,
  3.58,    3.58,    3.58,    3.58,
  3.61,    3.61,    3.61,    3.61,
  3.86,    3.86,    3.86,    3.86,
  3.3,     3.3,     3.3,     3.3,
  3.18,    3.18,    3.18,    3.18,
  2.67,    2.67,    2.67,    2.67,
  2.71,    2.71,    2.71,    2.71,
  2.87,    2.87,    2.87,    2.87,
  2.79,    2.79,    2.79,    2.79,
  2.51,    2.51,    2.51,    2.51,
  2.5,     2.5,     2.5,     2.5,
  2.65,    2.65,    2.65,    2.65,
  2.43,    2.43,    2.43,    2.43,
  2.24,    2.24,    2.24,    2.24,
  1.97,    1.97,    1.97,    1.97,
  2.2,     2.2,     2.2,     2.2,
  2.38,    2.38,    2.38,    2.38,
  2.39,    2.39,    2.39,    2.39,
  2.3,     2.3,     2.3,     2.3,
  2.53,    2.53,    2.53,    2.53,
  2.56,    2.56,    2.56,    2.56,
  2.46,    2.46,    2.46,    2.46,
  2.25,    2.25,    2.25,    2.25,
  2.11,    2.11,    2.11,    2.11,
  2.12,    2.12,    2.12,    2.12,
  2.21,    2.21,    2.21,    2.21,
  2.13,    2.13,    2.13,    2.13,
  1.84,    1.84,    1.84,    1.84,
  2.03,    2.03,    2.03,    2.03,
  2.68,    2.68,    2.68,    2.68,
  2.87,    2.87,    2.87,    2.87,
  3.18,    3.18,    3.18,    3.18,
  3.35,    3.35,    3.35,    3.35,
  2.59,    2.59,    2.59,    2.59,
  3.15,    3.15,    3.15,    3.15,
  2.87,    2.87,    2.87,    2.87,
  2.53,    2.53,    2.53,    2.53,
  2.81,    2.81,    2.81,    2.81,
  3.01,    3.01,    3.01,    3.01,
  2.27,    2.27,    2.27,    2.27,
  2.26,    2.26,    2.26,    2.26,
  2.31,    2.31,    2.31,    2.31,
  2.77,    2.77,    2.77,    2.77,
  3.12,    3.12,    3.12,    3.12,
  3.19,    3.19,    3.19,    3.19,
  3.23,    3.23,    3.23,    3.23,
  3.45,    3.45,    3.45,    3.45,
  3.06,    3.06,    3.06,    3.06,
  3.27,    3.27,    3.27,    3.27,
  2.99,    2.99,    2.99,    2.99,
  3.09,    3.09,    3.09,    3.09,
  2.81,    2.81,    2.81,    2.81,
  2.71,    2.71,    2.71,    2.71,
  2.26,    2.26,    2.26,    2.26,
  2.49,    2.49,    2.49,    2.49,
  2.36,    2.36,    2.36,    2.36,
  2.34,    2.34,    2.34,    2.34,
  2.31,    2.31,    2.31,    2.31,
  2.57,    2.57,    2.57,    2.57,
  2.67,    2.67,    2.67,    2.67,
  2.83,    2.83,    2.83,    2.83,
  3.11,    3.11,    3.11,    3.11,
  2.98,    2.98,    2.98,    2.98,
  2.79,    2.79,    2.79,    2.79,
  3.23,    3.23,    3.23,    3.23,
  3.08,    3.08,    3.08,    3.08,
  2.97,    2.97,    2.97,    2.97,
  3.09,    3.09,    3.09,    3.09,
  2.93,    2.93,    2.93,    2.93,
  3.1,     3.1,     3.1,     3.1,
  3.03,    3.03,    3.03,    3.03,
  3.05,    3.05,    3.05,    3.05,
  3.33,    3.33,    3.33,    3.33,
  3.05,    3.05,    3.05,    3.05,
  2.97,    2.97,    2.97,    2.97,
  2.63,    2.63,    2.63,    2.63,
  2.61,    2.61,    2.61,    2.61,
  2.54,    2.54,    2.54,    2.54,
  2.61,    2.61,    2.61,    2.61,
  2.44,    2.44,    2.44,    2.44,
  2.62,    2.62,    2.62,    2.62,
  3.17,    3.17,    3.17,    3.17,
  3.04,    3.04,    3.04,    3.04,
  2.84,    2.84,    2.84,    2.84,
  3.19,    3.19,    3.19,    3.19,
  3.32,    3.32,    3.32,    3.32,
  3.07,    3.07,    3.07,    3.07,
  3.29,    3.29,    3.29,    3.29,
  3.09,    3.09,    3.09,    3.09,
  3.16,    3.16,    3.16,    3.16,
  3.34,    3.34,    3.34,    3.34,
  2.94,    2.94,    2.94,    2.94,
  2.66,    2.66,    2.66,    2.66,
  2.71,    2.71,    2.71,    2.71,
  2.46,    2.46,    2.46,    2.46,
  2.37,    2.37,    2.37,    2.37,
  2.6,     2.6,     2.6,     2.6,
  2.52,    2.52,    2.52,    2.52,
  2.38,    2.38,    2.38,    2.38,
  2.59,    2.59,    2.59,    2.59,
  2.7,     2.7,     2.7,     2.7,
  2.87,    2.87,    2.87,    2.87,
  2.83,    2.83,    2.83,    2.83,
  3,       3,       3,       3,
  2.68,    2.68,    2.68,    2.68,
  2.7,     2.7,     2.7,     2.7,
  2.53,    2.53,    2.53,    2.53,
  2.63,    2.63,    2.63,    2.63,
  2.62,    2.62,    2.62,    2.62,
  2.48,    2.48,    2.48,    2.48,
  2.52,    2.52,    2.52,    2.52,
  2.47,    2.47,    2.47,    2.47,
  2.6,     2.6,     2.6,     2.6,
  2.64,    2.64,    2.64,    2.64,
  2.81,    2.81,    2.81,    2.81,
  2.64,    2.64,    2.64,    2.64,
  2.75,    2.75,    2.75,    2.75,
  2.45,    2.45,    2.45,    2.45,
  2.74,    2.74,    2.74,    2.74,
  2.64,    2.64,    2.64,    2.64,
  2.48,    2.48,    2.48,    2.48,
  2.52,    2.52,    2.52,    2.52,
  2.28,    2.28,    2.28,    2.28,
  2.17,    2.17,    2.17,    2.17,
  2.11,    2.11,    2.11,    2.11,
  2.22,    2.22,    2.22,    2.22,
  2.37,    2.37,    2.37,    2.37,
  2.41,    2.41,    2.41,    2.41,
  1.94,    1.94,    1.94,    1.94,
  2.08,    2.08,    2.08,    2.08,
  1.87,    1.87,    1.87,    1.87,
  1.48,    1.48,    1.48,    1.48,
  1.42,    1.42,    1.42,    1.42,
  0.97,    0.97,    0.97,    0.97,
  0.95,    0.95,    0.95,    0.95,
  1.08,    1.08,    1.08,    1.08,
  0.26,    0.26,    0.26,    0.26,
  0.53,    0.53,    0.53,    0.53,
  0.5,     0.5,     0.5,     0.5,
  0.98,    0.98,    0.98,    0.98,
  0.86,    0.86,    0.86,    0.86,
  1.15,    1.15,    1.15,    1.15,
  1.31,    1.31,    1.31,    1.31,
  1.63,    1.63,    1.63,    1.63,
  1.97,    1.97,    1.97,    1.97,
  1.77,    1.77,    1.77,    1.77,
  2.07,    2.07,    2.07,    2.07,
  3.05,    3.05,    3.05,    3.05,
  4.64,    4.64,    4.64,    4.64,
  4.92,    4.92,    4.92,    4.92,
  4.28,    4.28,    4.28,    4.28,
  3.79,    3.79,    3.79,    3.79,
  2.95,    2.95,    2.95,    2.95,
  2.47,    2.47,    2.47,    2.47,
  2.07,    2.07,    2.07,    2.07,
  2.16,    2.16,    2.16,    2.16,
  2.58,    2.58,    2.58,    2.58,
  1.85,    1.85,    1.85,    1.85,
  2.15,    2.15,    2.15,    2.15,
  1.69,    1.69,    1.69,    1.69,
  2.36,    2.36,    2.36,    2.36,
  2.11,    2.11,    2.11,    2.11,
  2.01,    2.01,    2.01,    2.01,
  2.07,    2.07,    2.07,    2.07,
  2.36,    2.36,    2.36,    2.36,
  2.21,    2.21,    2.21,    2.21,
  2.16,    2.16,    2.16,    2.16,
  2.52,    2.52,    2.52,    2.52,
  1.6,     1.6,     1.6,     1.6,
  0.41,    0.41,    0.41,    0.41,
  1.37,    1.37,    1.37,    1.37,
  1.67,    1.67,    1.67,    1.67,
  1.91,    1.91,    1.91,    1.91,
  1.92,    1.92,    1.92,    1.92,
  1.79,    1.79,    1.79,    1.79,
  1.87,    1.87,    1.87,    1.87,
  1.99,    1.99,    1.99,    1.99,
  1.66,    1.66,    1.66,    1.66,
  2.16,    2.16,    2.16,    2.16,
  1.16,    1.16,    1.16,    1.16,
  1.15,    1.15,    1.15,    1.15,
  1.5,     1.5,     1.5,     1.5,
  2.18,    2.18,    2.18,    2.18,
  1.71,    1.71,    1.71,    1.71,
  1.38,    1.38,    1.38,    1.38,
  1.95,    1.95,    1.95,    1.95,
  1.48,    1.48,    1.48,    1.48,
  1.4,     1.4,     1.4,     1.4,
  1.67,    1.67,    1.67,    1.67,
  2.03,    2.03,    2.03,    2.03,
  1.79,    1.79,    1.79,    1.79,
  1.88,    1.88,    1.88,    1.88,
  1.79,    1.79,    1.79,    1.79,
  1.89,    1.89,    1.89,    1.89,
  2.13,    2.13,    2.13,    2.13,
  2.02,    2.02,    2.02,    2.02,
  2.04,    2.04,    2.04,    2.04,
  2.05,    2.05,    2.05,    2.05,
  1.7,     1.7,     1.7,     1.7,
  2.04,    2.04,    2.04,    2.04,
  2.25,    2.25,    2.25,    2.25,
  1.87,    1.87,    1.87,    1.87,
  1.63,    1.63,    1.63,    1.63,
  1.96,    1.96,    1.96,    1.96,
  2.1,     2.1,     2.1,     2.1,
  2.13,    2.13,    2.13,    2.13,
  1.99,    1.99,    1.99,    1.99,
  1.59,    1.59,    1.59,    1.59,
  1.55,    1.55,    1.55,    1.55,
  2.01,    2.01,    2.01,    2.01,
  1.94,    1.94,    1.94,    1.94,
  2.11,    2.11,    2.11,    2.11,
  2.19,    2.19,    2.19,    2.19,
  1.9,     1.9,     1.9,     1.9,
  1.59,    1.59,    1.59,    1.59,
  1.97,    1.97,    1.97,    1.97,
  1.72,    1.72,    1.72,    1.72,
  1.94,    1.94,    1.94,    1.94,
  2.09,    2.09,    2.09,    2.09,
  2.26,    2.26,    2.26,    2.26,
  2.28,    2.28,    2.28,    2.28,
  2.56,    2.56,    2.56,    2.56,
  2.55,    2.55,    2.55,    2.55,
  2.33,    2.33,    2.33,    2.33,
  1.9,     1.9,     1.9,     1.9,
  2.17,    2.17,    2.17,    2.17,
  2.37,    2.37,    2.37,    2.37,
  2.43,    2.43,    2.43,    2.43,
  2.49,    2.49,    2.49,    2.49,
  2.72,    2.72,    2.72,    2.72,
  3.02,    3.02,    3.02,    3.02,
  2.79,    2.79,    2.79,    2.79,
  3.01,    3.01,    3.01,    3.01,
  2.95,    2.95,    2.95,    2.95,
  2.76,    2.76,    2.76,    2.76,
  2.5,     2.5,     2.5,     2.5,
  2.24,    2.24,    2.24,    2.24,
  2.77,    2.77,    2.77,    2.77,
  3.14,    3.14,    3.14,    3.14,
  3.27,    3.27,    3.27,    3.27,
  3.18,    3.18,    3.18,    3.18,
  3.15,    3.15,    3.15,    3.15,
  3.3,     3.3,     3.3,     3.3,
  2.67,    2.67,    2.67,    2.67,
  2.81,    2.81,    2.81,    2.81,
  2.95,    2.95,    2.95,    2.95,
  2.83,    2.83,    2.83,    2.83,
  2.46,    2.46,    2.46,    2.46,
  2.5,     2.5,     2.5,     2.5,
  2.51,    2.51,    2.51,    2.51,
  2.3,     2.3,     2.3,     2.3,
  2.62,    2.62,    2.62,    2.62,
  2.92,    2.92,    2.92,    2.92,
  3.01,    3.01,    3.01,    3.01,
  2.53,    2.53,    2.53,    2.53,
  2.84,    2.84,    2.84,    2.84,
  3.72,    3.72,    3.72,    3.72,
  3.1,     3.1,     3.1,     3.1,
  2.97,    2.97,    2.97,    2.97,
  2.9,     2.9,     2.9,     2.9,
  2.74,    2.74,    2.74,    2.74,
  2.35,    2.35,    2.35,    2.35,
  2.07,    2.07,    2.07,    2.07,
  2.01,    2.01,    2.01,    2.01,
  2.01,    2.01,    2.01,    2.01,
  1.97,    1.97,    1.97,    1.97,
  2.21,    2.21,    2.21,    2.21,
  1.98,    1.98,    1.98,    1.98,
  1.88,    1.88,    1.88,    1.88,
  1.7,     1.7,     1.7,     1.7,
  1.32,    1.32,    1.32,    1.32,
  1.17,    1.17,    1.17,    1.17,
  1.49,    1.49,    1.49,    1.49,
  1.61,    1.61,    1.61,    1.61,
  1.31,    1.31,    1.31,    1.31,
  1.38,    1.38,    1.38,    1.38,
  1.58,    1.58,    1.58,    1.58,
  1.65,    1.65,    1.65,    1.65,
  2.34,    2.34,    2.34,    2.34,
  2.71,    2.71,    2.71,    2.71,
  2.66,    2.66,    2.66,    2.66,
  2.76,    2.76,    2.76,    2.76,
  3.2,     3.2,     3.2,     3.2,
  2.3,     2.3,     2.3,     2.3,
  2.29,    2.29,    2.29,    2.29,
  2.06,    2.06,    2.06,    2.06,
  1.68,    1.68,    1.68,    1.68,
  1.65,    1.65,    1.65,    1.65,
  1.87,    1.87,    1.87,    1.87,
  2.49,    2.49,    2.49,    2.49,
  2.46,    2.46,    2.46,    2.46,
  2.73,    2.73,    2.73,    2.73,
  1.99,    1.99,    1.99,    1.99,
  1.73,    1.73,    1.73,    1.73,
  1.66,    1.66,    1.66,    1.66,
  1.77,    1.77,    1.77,    1.77,
  1.76,    1.76,    1.76,    1.76,
  1.64,    1.64,    1.64,    1.64,
  1.67,    1.67,    1.67,    1.67,
  1.56,    1.56,    1.56,    1.56,
  1.63,    1.63,    1.63,    1.63,
  1.73,    1.73,    1.73,    1.73,
  1.55,    1.55,    1.55,    1.55,
  1.82,    1.82,    1.82,    1.82,
  1.89,    1.89,    1.89,    1.89,
  1.79,    1.79,    1.79,    1.79,
  1.84,    1.84,    1.84,    1.84,
  1.67,    1.67,    1.67,    1.67,
  1.39,    1.39,    1.39,    1.39,
  1.37,    1.37,    1.37,    1.37,
  1.33,    1.33,    1.33,    1.33,
  1.48,    1.48,    1.48,    1.48,
  1.53,    1.53,    1.53,    1.53,
  1.69,    1.69,    1.69,    1.69,
  1.6,     1.6,     1.6,     1.6,
  1.57,    1.57,    1.57,    1.57,
  1.98,    1.98,    1.98,    1.98,
  1.82,    1.82,    1.82,    1.82,
  2.04,    2.04,    2.04,    2.04,
  1.84,    1.84,    1.84,    1.84,
  1.46,    1.46,    1.46,    1.46,
  2.29,    2.29,    2.29,    2.29,
  2.25,    2.25,    2.25,    2.25,
  1.85,    1.85,    1.85,    1.85,
  1.65,    1.65,    1.65,    1.65,
  1.71,    1.71,    1.71,    1.71,
  1.79,    1.79,    1.79,    1.79,
  1.59,    1.59,    1.59,    1.59,
  1.55,    1.55,    1.55,    1.55,
  2.09,    2.09,    2.09,    2.09,
  1.89,    1.89,    1.89,    1.89,
  1.97,    1.97,    1.97,    1.97,
  1.43,    1.43,    1.43,    1.43,
  1.22,    1.22,    1.22,    1.22,
  0.69,    0.69,    0.69,    0.69,
  2.07,    2.07,    2.07,    2.07,
  1.99,    1.99,    1.99,    1.99,
  1.94,    1.94,    1.94,    1.94,
  0.88,    0.88,    0.88,    0.88,
  0.59,    0.59,    0.59,    0.59,
  1.58,    1.58,    1.58,    1.58,
  1.18,    1.18,    1.18,    1.18,
  0.75,    0.75,    0.75,    0.75,
  0.54,    0.54,    0.54,    0.54,
  1.23,    1.23,    1.23,    1.23,
  1.46,    1.46,    1.46,    1.46,
  1.13,    1.13,    1.13,    1.13,
  1.25,    1.25,    1.25,    1.25,
  1.44,    1.44,    1.44,    1.44,
  1.58,    1.58,    1.58,    1.58,
  1.64,    1.64,    1.64,    1.64,
  1.31,    1.31,    1.31,    1.31,
  1.69,    1.69,    1.69,    1.69,
  1.7,     1.7,     1.7,     1.7,
  1.82,    1.82,    1.82,    1.82,
  1.36,    1.36,    1.36,    1.36,
  1.26,    1.26,    1.26,    1.26,
  1.89,    1.89,    1.89,    1.89,
  1.79,    1.79,    1.79,    1.79,
  1.7,     1.7,     1.7,     1.7,
  1.31,    1.31,    1.31,    1.31,
  1.95,    1.95,    1.95,    1.95,
  1.72,    1.72,    1.72,    1.72,
  1.75,    1.75,    1.75,    1.75,
  1.9,     1.9,     1.9,     1.9,
  1.86,    1.86,    1.86,    1.86,
  1.86,    1.86,    1.86,    1.86,
  1.62,    1.62,    1.62,    1.62,
  1.03,    1.03,    1.03,    1.03,
  1.72,    1.72,    1.72,    1.72,
  2.33,    2.33,    2.33,    2.33,
  2.02,    2.02,    2.02,    2.02,
  2.02,    2.02,    2.02,    2.02,
  2.33,    2.33,    2.33,    2.33,
  2.35,    2.35,    2.35,    2.35,
  2.68,    2.68,    2.68,    2.68,
  2.24,    2.24,    2.24,    2.24,
  2.53,    2.53,    2.53,    2.53,
  2.33,    2.33,    2.33,    2.33,
  2.33,    2.33,    2.33,    2.33,
  2.15,    2.15,    2.15,    2.15,
  2.63,    2.63,    2.63,    2.63,
  2.46,    2.46,    2.46,    2.46,
  2.25,    2.25,    2.25,    2.25,
  2.09,    2.09,    2.09,    2.09,
  1.91,    1.91,    1.91,    1.91,
  1.8,     1.8,     1.8,     1.8,
  1.96,    1.96,    1.96,    1.96,
  2.21,    2.21,    2.21,    2.21,
  2.2,     2.2,     2.2,     2.2,
  2.17,    2.17,    2.17,    2.17,
  2.09,    2.09,    2.09,    2.09,
  2.29,    2.29,    2.29,    2.29,
  2.52,    2.52,    2.52,    2.52,
  2.38,    2.38,    2.38,    2.38,
  2.5,     2.5,     2.5,     2.5,
  2.65,    2.65,    2.65,    2.65,
  2.75,    2.75,    2.75,    2.75,
  2.57,    2.57,    2.57,    2.57,
  2.95,    2.95,    2.95,    2.95,
  3.33,    3.33,    3.33,    3.33,
  3.01,    3.01,    3.01,    3.01,
  2.96,    2.96,    2.96,    2.96,
  3.39,    3.39,    3.39,    3.39,
  3.33,    3.33,    3.33,    3.33,
  3.23,    3.23,    3.23,    3.23,
  3.39,    3.39,    3.39,    3.39,
  3.26,    3.26,    3.26,    3.26,
  3.56,    3.56,    3.56,    3.56,
  3.8,     3.8,     3.8,     3.8,
  3.71,    3.71,    3.71,    3.71,
  3.93,    3.93,    3.93,    3.93,
  4.28,    4.28,    4.28,    4.28,
  4.4,     4.4,     4.4,     4.4,
  4.6,     4.6,     4.6,     4.6,
  4.61,    4.61,    4.61,    4.61,
  4.07,    4.07,    4.07,    4.07,
  3.9,     3.9,     3.9,     3.9,
  4.26,    4.26,    4.26,    4.26,
  3.74,    3.74,    3.74,    3.74,
  4.31,    4.31,    4.31,    4.31,
  4.27,    4.27,    4.27,    4.27,
  4.24,    4.24,    4.24,    4.24,
  4.57,    4.57,    4.57,    4.57,
  4.49,    4.49,    4.49,    4.49,
  4.35,    4.35,    4.35,    4.35,
  4.42,    4.42,    4.42,    4.42,
  4.02,    4.02,    4.02,    4.02,
  3.7,     3.7,     3.7,     3.7,
  3.58,    3.58,    3.58,    3.58,
  3.47,    3.47,    3.47,    3.47,
  3.13,    3.13,    3.13,    3.13,
  2.99,    2.99,    2.99,    2.99,
  3.45,    3.45,    3.45,    3.45,
  3.6,     3.6,     3.6,     3.6,
  4,       4,       4,       4,
  3.77,    3.77,    3.77,    3.77,
  3.95,    3.95,    3.95,    3.95,
  4.09,    4.09,    4.09,    4.09,
  3.78,    3.78,    3.78,    3.78,
  4.02,    4.02,    4.02,    4.02,
  4.16,    4.16,    4.16,    4.16,
  3.98,    3.98,    3.98,    3.98,
  3.48,    3.48,    3.48,    3.48,
  3.32,    3.32,    3.32,    3.32,
  3.64,    3.64,    3.64,    3.64,
  3.43,    3.43,    3.43,    3.43,
  3.42,    3.42,    3.42,    3.42,
  3.87,    3.87,    3.87,    3.87,
  3.34,    3.34,    3.34,    3.34,
  3.51,    3.51,    3.51,    3.51,
  3.23,    3.23,    3.23,    3.23,
  3.31,    3.31,    3.31,    3.31,
  2.8,     2.8,     2.8,     2.8,
  1.98,    1.98,    1.98,    1.98,
  2.02,    2.02,    2.02,    2.02,
  2.22,    2.22,    2.22,    2.22,
  2.25,    2.25,    2.25,    2.25,
  2.44,    2.44,    2.44,    2.44,
  2.04,    2.04,    2.04,    2.04,
  2.22,    2.22,    2.22,    2.22,
  2.5,     2.5,     2.5,     2.5,
  2.78,    2.78,    2.78,    2.78,
  2.73,    2.73,    2.73,    2.73,
  3.1,     3.1,     3.1,     3.1,
  2.99,    2.99,    2.99,    2.99,
  2.97,    2.97,    2.97,    2.97,
  3.11,    3.11,    3.11,    3.11,
  2.85,    2.85,    2.85,    2.85,
  2.98,    2.98,    2.98,    2.98,
  2.83,    2.83,    2.83,    2.83,
  3.08,    3.08,    3.08,    3.08,
  2.72,    2.72,    2.72,    2.72,
  2.65,    2.65,    2.65,    2.65,
  2.18,    2.18,    2.18,    2.18,
  2.14,    2.14,    2.14,    2.14,
  2.45,    2.45,    2.45,    2.45,
  2.61,    2.61,    2.61,    2.61,
  2.45,    2.45,    2.45,    2.45,
  2.52,    2.52,    2.52,    2.52,
  2.82,    2.82,    2.82,    2.82,
  3.13,    3.13,    3.13,    3.13,
  2.94,    2.94,    2.94,    2.94,
  3.01,    3.01,    3.01,    3.01,
  2.85,    2.85,    2.85,    2.85,
  2.85,    2.85,    2.85,    2.85,
  2.46,    2.46,    2.46,    2.46,
  2.59,    2.59,    2.59,    2.59,
  2.43,    2.43,    2.43,    2.43,
  2.43,    2.43,    2.43,    2.43,
  2.41,    2.41,    2.41,    2.41,
  2.51,    2.51,    2.51,    2.51,
  3.16,    3.16,    3.16,    3.16,
  2.96,    2.96,    2.96,    2.96,
  3.49,    3.49,    3.49,    3.49,
  3.64,    3.64,    3.64,    3.64,
  3.81,    3.81,    3.81,    3.81,
  4.22,    4.22,    4.22,    4.22,
  3.92,    3.92,    3.92,    3.92,
  4.08,    4.08,    4.08,    4.08,
  4.45,    4.45,    4.45,    4.45,
  4.29,    4.29,    4.29,    4.29,
  4.09,    4.09,    4.09,    4.09,
  3.67,    3.67,    3.67,    3.67,
  3.44,    3.44,    3.44,    3.44,
  3.19,    3.19,    3.19,    3.19,
  3.25,    3.25,    3.25,    3.25,
  3.4,     3.4,     3.4,     3.4,
  3.37,    3.37,    3.37,    3.37,
  3.48,    3.48,    3.48,    3.48,
  3.52,    3.52,    3.52,    3.52,
  2.95,    2.95,    2.95,    2.95,
  3.35,    3.35,    3.35,    3.35,
  3.58,    3.58,    3.58,    3.58,
  3.44,    3.44,    3.44,    3.44,
  3.31,    3.31,    3.31,    3.31,
  3.91,    3.91,    3.91,    3.91,
  4.4,     4.4,     4.4,     4.4,
  4.21,    4.21,    4.21,    4.21,
  4.67,    4.67,    4.67,    4.67,
  4.68,    4.68,    4.68,    4.68,
  4.59,    4.59,    4.59,    4.59,
  4.15,    4.15,    4.15,    4.15,
  3.79,    3.79,    3.79,    3.79,
  3.88,    3.88,    3.88,    3.88,
  3.87,    3.87,    3.87,    3.87,
  3.89,    3.89,    3.89,    3.89,
  4.01,    4.01,    4.01,    4.01,
  4.12,    4.12,    4.12,    4.12,
  3.64,    3.64,    3.64,    3.64,
  3.62,    3.62,    3.62,    3.62,
  3.18,    3.18,    3.18,    3.18,
  2.96,    2.96,    2.96,    2.96,
  3.15,    3.15,    3.15,    3.15,
  2.93,    2.93,    2.93,    2.93,
  3.47,    3.47,    3.47,    3.47,
  3.66,    3.66,    3.66,    3.66,
  3.18,    3.18,    3.18,    3.18,
  3.23,    3.23,    3.23,    3.23,
  3.08,    3.08,    3.08,    3.08,
  3.47,    3.47,    3.47,    3.47,
  3.3,     3.3,     3.3,     3.3,
  3.49,    3.49,    3.49,    3.49,
  3.85,    3.85,    3.85,    3.85,
  3.47,    3.47,    3.47,    3.47,
  3.08,    3.08,    3.08,    3.08,
  3.78,    3.78,    3.78,    3.78,
  3.66,    3.66,    3.66,    3.66,
  3.31,    3.31,    3.31,    3.31,
  3.43,    3.43,    3.43,    3.43,
  3.79,    3.79,    3.79,    3.79,
  3.45,    3.45,    3.45,    3.45,
  3.62,    3.62,    3.62,    3.62,
  3.56,    3.56,    3.56,    3.56,
  3.42,    3.42,    3.42,    3.42,
  3.27,    3.27,    3.27,    3.27,
  3.4,     3.4,     3.4,     3.4,
  3.17,    3.17,    3.17,    3.17,
  2.99,    2.99,    2.99,    2.99,
  3.6,     3.6,     3.6,     3.6,
  3.99,    3.99,    3.99,    3.99,
  3.7,     3.7,     3.7,     3.7,
  3.9,     3.9,     3.9,     3.9,
  3.39,    3.39,    3.39,    3.39,
  3.94,    3.94,    3.94,    3.94,
  4.05,    4.05,    4.05,    4.05,
  3.92,    3.92,    3.92,    3.92,
  3.91,    3.91,    3.91,    3.91,
  3.8,     3.8,     3.8,     3.8,
  3.4,     3.4,     3.4,     3.4,
  3.67,    3.67,    3.67,    3.67,
  3.53,    3.53,    3.53,    3.53,
  3.89,    3.89,    3.89,    3.89,
  3.77,    3.77,    3.77,    3.77,
  3.72,    3.72,    3.72,    3.72,
  4.11,    4.11,    4.11,    4.11,
  3.92,    3.92,    3.92,    3.92,
  4.2,     4.2,     4.2,     4.2,
  4.29,    4.29,    4.29,    4.29,
  3.66,    3.66,    3.66,    3.66,
  4.23,    4.23,    4.23,    4.23,
  4.41,    4.41,    4.41,    4.41,
  3.97,    3.97,    3.97,    3.97,
  4.08,    4.08,    4.08,    4.08,
  3.99,    3.99,    3.99,    3.99,
  3.97,    3.97,    3.97,    3.97,
  4.03,    4.03,    4.03,    4.03,
  3.77,    3.77,    3.77,    3.77,
  4.19,    4.19,    4.19,    4.19,
  4.38,    4.38,    4.38,    4.38,
  4.09,    4.09,    4.09,    4.09,
  5.19,    5.19,    5.19,    5.19,
  4.52,    4.52,    4.52,    4.52,
  4.03,    4.03,    4.03,    4.03,
  4.02,    4.02,    4.02,    4.02,
  4.43,    4.43,    4.43,    4.43,
  4.58,    4.58,    4.58,    4.58,
  4.55,    4.55,    4.55,    4.55,
  5.24,    5.24,    5.24,    5.24,
  5.16,    5.16,    5.16,    5.16,
  4.29,    4.29,    4.29,    4.29,
  4.49,    4.49,    4.49,    4.49,
  4.76,    4.76,    4.76,    4.76,
  4.43,    4.43,    4.43,    4.43,
  4.53,    4.53,    4.53,    4.53,
  4.92,    4.92,    4.92,    4.92,
  5.54,    5.54,    5.54,    5.54,
  4.57,    4.57,    4.57,    4.57,
  5.78,    5.78,    5.78,    5.78,
  5.82,    5.82,    5.82,    5.82,
  5.77,    5.77,    5.77,    5.77,
  5.94,    5.94,    5.94,    5.94,
  5.44,    5.44,    5.44,    5.44,
  5.6,     5.6,     5.6,     5.6,
  5.74,    5.74,    5.74,    5.74,
  5.02,    5.02,    5.02,    5.02,
  4.75,    4.75,    4.75,    4.75,
  4.17,    4.17,    4.17,    4.17,
  4.2,     4.2,     4.2,     4.2,
  4.6,     4.6,     4.6,     4.6,
  5.23,    5.23,    5.23,    5.23,
  4.47,    4.47,    4.47,    4.47,
  4.78,    4.78,    4.78,    4.78,
  5.44,    5.44,    5.44,    5.44,
  5.16,    5.16,    5.16,    5.16,
  5.25,    5.25,    5.25,    5.25,
  4.96,    4.96,    4.96,    4.96,
  4.86,    4.86,    4.86,    4.86,
  5.03,    5.03,    5.03,    5.03,
  4.73,    4.73,    4.73,    4.73,
  5.52,    5.52,    5.52,    5.52,
  5.77,    5.77,    5.77,    5.77,
  5.66,    5.66,    5.66,    5.66,
  5.47,    5.47,    5.47,    5.47,
  5.04,    5.04,    5.04,    5.04,
  5.94,    5.94,    5.94,    5.94,
  4.76,    4.76,    4.76,    4.76,
  4.47,    4.47,    4.47,    4.47,
  4.16,    4.16,    4.16,    4.16,
  4.23,    4.23,    4.23,    4.23,
  4.3,     4.3,     4.3,     4.3,
  3.99,    3.99,    3.99,    3.99,
  3.11,    3.11,    3.11,    3.11,
  2.91,    2.91,    2.91,    2.91,
  3.11,    3.11,    3.11,    3.11,
  2.89,    2.89,    2.89,    2.89,
  2.59,    2.59,    2.59,    2.59,
  2.75,    2.75,    2.75,    2.75,
  2.66,    2.66,    2.66,    2.66,
  2.79,    2.79,    2.79,    2.79,
  2.87,    2.87,    2.87,    2.87,
  3.02,    3.02,    3.02,    3.02,
  3.21,    3.21,    3.21,    3.21,
  3.39,    3.39,    3.39,    3.39,
  3.21,    3.21,    3.21,    3.21,
  3.14,    3.14,    3.14,    3.14,
  3.85,    3.85,    3.85,    3.85,
  4.17,    4.17,    4.17,    4.17,
  4.5,     4.5,     4.5,     4.5,
  3.86,    3.86,    3.86,    3.86,
  4.13,    4.13,    4.13,    4.13,
  4.69,    4.69,    4.69,    4.69,
  4.77,    4.77,    4.77,    4.77,
  4.47,    4.47,    4.47,    4.47,
  5.22,    5.22,    5.22,    5.22,
  4.16,    4.16,    4.16,    4.16,
  4.4,     4.4,     4.4,     4.4,
  3.96,    3.96,    3.96,    3.96,
  4.34,    4.34,    4.34,    4.34,
  4.28,    4.28,    4.28,    4.28,
  3.94,    3.94,    3.94,    3.94,
  4.01,    4.01,    4.01,    4.01,
  3.43,    3.43,    3.43,    3.43,
  4.32,    4.32,    4.32,    4.32,
  3.76,    3.76,    3.76,    3.76,
  3.39,    3.39,    3.39,    3.39,
  3.25,    3.25,    3.25,    3.25,
  3.55,    3.55,    3.55,    3.55,
  3.46,    3.46,    3.46,    3.46,
  4,       4,       4,       4,
  3.83,    3.83,    3.83,    3.83,
  3.16,    3.16,    3.16,    3.16,
  3.47,    3.47,    3.47,    3.47,
  3.52,    3.52,    3.52,    3.52,
  3.24,    3.24,    3.24,    3.24,
  3.1,     3.1,     3.1,     3.1,
  2.68,    2.68,    2.68,    2.68,
  2.91,    2.91,    2.91,    2.91,
  2.52,    2.52,    2.52,    2.52,
  2.68,    2.68,    2.68,    2.68,
  2.69,    2.69,    2.69,    2.69,
  4.28,    4.28,    4.28,    4.28,
  4.92,    4.92,    4.92,    4.92,
  3.81,    3.81,    3.81,    3.81,
  3.21,    3.21,    3.21,    3.21,
  2.97,    2.97,    2.97,    2.97,
  3.56,    3.56,    3.56,    3.56,
  3.69,    3.69,    3.69,    3.69,
  3.9,     3.9,     3.9,     3.9,
  3.84,    3.84,    3.84,    3.84,
  3.31,    3.31,    3.31,    3.31,
  5.04,    5.04,    5.04,    5.04,
  4.85,    4.85,    4.85,    4.85,
  3.31,    3.31,    3.31,    3.31,
  2.93,    2.93,    2.93,    2.93,
  3.38,    3.38,    3.38,    3.38,
  3.43,    3.43,    3.43,    3.43,
  3.51,    3.51,    3.51,    3.51,
  3.65,    3.65,    3.65,    3.65,
  3.69,    3.69,    3.69,    3.69,
  3.68,    3.68,    3.68,    3.68,
  4.12,    4.12,    4.12,    4.12,
  3.31,    3.31,    3.31,    3.31,
  3.42,    3.42,    3.42,    3.42,
  3.51,    3.51,    3.51,    3.51,
  3.4,     3.4,     3.4,     3.4,
  3.83,    3.83,    3.83,    3.83,
  3.6,     3.6,     3.6,     3.6,
  3.94,    3.94,    3.94,    3.94,
  4.15,    4.15,    4.15,    4.15,
  4.5,     4.5,     4.5,     4.5,
  4.14,    4.14,    4.14,    4.14,
  3.62,    3.62,    3.62,    3.62,
  3.75,    3.75,    3.75,    3.75,
  3.58,    3.58,    3.58,    3.58,
  3.36,    3.36,    3.36,    3.36,
  3.34,    3.34,    3.34,    3.34,
  3.53,    3.53,    3.53,    3.53,
  2.97,    2.97,    2.97,    2.97,
  3.28,    3.28,    3.28,    3.28,
  3.54,    3.54,    3.54,    3.54,
  3.49,    3.49,    3.49,    3.49,
  3.32,    3.32,    3.32,    3.32,
  2.81,    2.81,    2.81,    2.81,
  2.77,    2.77,    2.77,    2.77,
  2.91,    2.91,    2.91,    2.91,
  2.44,    2.44,    2.44,    2.44,
  2.34,    2.34,    2.34,    2.34,
  2.55,    2.55,    2.55,    2.55,
  2.65,    2.65,    2.65,    2.65,
  2.37,    2.37,    2.37,    2.37,
  2.2,     2.2,     2.2,     2.2,
  2.22,    2.22,    2.22,    2.22,
  2.11,    2.11,    2.11,    2.11,
  2.08,    2.08,    2.08,    2.08,
  2.27,    2.27,    2.27,    2.27,
  2.22,    2.22,    2.22,    2.22,
  2.31,    2.31,    2.31,    2.31,
  2.42,    2.42,    2.42,    2.42,
  2.13,    2.13,    2.13,    2.13,
  1.65,    1.65,    1.65,    1.65,
  1.62,    1.62,    1.62,    1.62,
  1.45,    1.45,    1.45,    1.45,
  1.92,    1.92,    1.92,    1.92,
  1.91,    1.91,    1.91,    1.91,
  1.83,    1.83,    1.83,    1.83,
  2.64,    2.64,    2.64,    2.64,
  3.33,    3.33,    3.33,    3.33,
  3.32,    3.32,    3.32,    3.32,
  3.14,    3.14,    3.14,    3.14,
  2.76,    2.76,    2.76,    2.76,
  2.47,    2.47,    2.47,    2.47,
  1.83,    1.83,    1.83,    1.83,
  2.16,    2.16,    2.16,    2.16,
  2.06,    2.06,    2.06,    2.06,
  2.8,     2.8,     2.8,     2.8,
  2.49,    2.49,    2.49,    2.49,
  3.3,     3.3,     3.3,     3.3,
  2.99,    2.99,    2.99,    2.99,
  3.54,    3.54,    3.54,    3.54,
  3.11,    3.11,    3.11,    3.11,
  2.87,    2.87,    2.87,    2.87,
  2.52,    2.52,    2.52,    2.52,
  2.17,    2.17,    2.17,    2.17,
  2.11,    2.11,    2.11,    2.11,
  2.24,    2.24,    2.24,    2.24,
  2.08,    2.08,    2.08,    2.08,
  1.98,    1.98,    1.98,    1.98,
  1.9,     1.9,     1.9,     1.9,
  1.9,     1.9,     1.9,     1.9,
  1.72,    1.72,    1.72,    1.72,
  1.61,    1.61,    1.61,    1.61,
  1.56,    1.56,    1.56,    1.56,
  1.38,    1.38,    1.38,    1.38,
  1.96,    1.96,    1.96,    1.96,
  1.97,    1.97,    1.97,    1.97,
  2.26,    2.26,    2.26,    2.26,
  2.11,    2.11,    2.11,    2.11,
  2.21,    2.21,    2.21,    2.21,
  2.54,    2.54,    2.54,    2.54,
  2.19,    2.19,    2.19,    2.19,
  1.61,    1.61,    1.61,    1.61,
  2.09,    2.09,    2.09,    2.09,
  1.56,    1.56,    1.56,    1.56,
  2.16,    2.16,    2.16,    2.16,
  1.9,     1.9,     1.9,     1.9,
  1.98,    1.98,    1.98,    1.98,
  1.78,    1.78,    1.78,    1.78,
  2.24,    2.24,    2.24,    2.24,
  1.68,    1.68,    1.68,    1.68,
  1.37,    1.37,    1.37,    1.37,
  1.93,    1.93,    1.93,    1.93,
  2.28,    2.28,    2.28,    2.28,
  2.64,    2.64,    2.64,    2.64,
  3.43,    3.43,    3.43,    3.43,
  2.71,    2.71,    2.71,    2.71,
  3.14,    3.14,    3.14,    3.14,
  3.8,     3.8,     3.8,     3.8,
  3.28,    3.28,    3.28,    3.28,
  3.46,    3.46,    3.46,    3.46,
  2.43,    2.43,    2.43,    2.43,
  3.07,    3.07,    3.07,    3.07,
  2.77,    2.77,    2.77,    2.77,
  2.45,    2.45,    2.45,    2.45,
  3.33,    3.33,    3.33,    3.33,
  3,       3,       3,       3,
  3.54,    3.54,    3.54,    3.54,
  3.66,    3.66,    3.66,    3.66,
  4.11,    4.11,    4.11,    4.11,
  3.81,    3.81,    3.81,    3.81,
  3.84,    3.84,    3.84,    3.84,
  3.55,    3.55,    3.55,    3.55,
  3.62,    3.62,    3.62,    3.62,
  3.89,    3.89,    3.89,    3.89,
  4.02,    4.02,    4.02,    4.02,
  4.05,    4.05,    4.05,    4.05,
  3.79,    3.79,    3.79,    3.79,
  3.68,    3.68,    3.68,    3.68,
  3.16,    3.16,    3.16,    3.16,
  3.13,    3.13,    3.13,    3.13,
  3.58,    3.58,    3.58,    3.58,
  3.35,    3.35,    3.35,    3.35,
  2.55,    2.55,    2.55,    2.55,
  2.41,    2.41,    2.41,    2.41,
  2.67,    2.67,    2.67,    2.67,
  2.28,    2.28,    2.28,    2.28,
  2.48,    2.48,    2.48,    2.48,
  2.57,    2.57,    2.57,    2.57,
  2.67,    2.67,    2.67,    2.67,
  3.01,    3.01,    3.01,    3.01,
  3.79,    3.79,    3.79,    3.79,
  3.74,    3.74,    3.74,    3.74,
  4.08,    4.08,    4.08,    4.08,
  4.01,    4.01,    4.01,    4.01,
  4.48,    4.48,    4.48,    4.48,
  4.65,    4.65,    4.65,    4.65,
  3.74,    3.74,    3.74,    3.74,
  3.66,    3.66,    3.66,    3.66,
  4.3,     4.3,     4.3,     4.3,
  4.75,    4.75,    4.75,    4.75,
  4.15,    4.15,    4.15,    4.15,
  4.45,    4.45,    4.45,    4.45,
  4.14,    4.14,    4.14,    4.14,
  4.28,    4.28,    4.28,    4.28,
  4.61,    4.61,    4.61,    4.61,
  6.13,    6.13,    6.13,    6.13,
  6,       6,       6,       6,
  5.5,     5.5,     5.5,     5.5,
  5.41,    5.41,    5.41,    5.41,
  5.97,    5.97,    5.97,    5.97,
  5.87,    5.87,    5.87,    5.87,
  5.4,     5.4,     5.4,     5.4,
  5.45,    5.45,    5.45,    5.45,
  4.94,    4.94,    4.94,    4.94,
  5.44,    5.44,    5.44,    5.44,
  5.5,     5.5,     5.5,     5.5,
  5.53,    5.53,    5.53,    5.53,
  5.99,    5.99,    5.99,    5.99,
  5.07,    5.07,    5.07,    5.07,
  4.29,    4.29,    4.29,    4.29,
  4.39,    4.39,    4.39,    4.39,
  4.59,    4.59,    4.59,    4.59,
  4.05,    4.05,    4.05,    4.05,
  3.72,    3.72,    3.72,    3.72,
  4.02,    4.02,    4.02,    4.02,
  3.85,    3.85,    3.85,    3.85,
  3.8,     3.8,     3.8,     3.8,
  3.72,    3.72,    3.72,    3.72,
  4.13,    4.13,    4.13,    4.13,
  4.32,    4.32,    4.32,    4.32,
  4.25,    4.25,    4.25,    4.25,
  4.33,    4.33,    4.33,    4.33,
  4.35,    4.35,    4.35,    4.35,
  4.43,    4.43,    4.43,    4.43,
  5.11,    5.11,    5.11,    5.11,
  5.06,    5.06,    5.06,    5.06,
  4.98,    4.98,    4.98,    4.98,
  5.71,    5.71,    5.71,    5.71,
  5.41,    5.41,    5.41,    5.41,
  5.49,    5.49,    5.49,    5.49,
  5.7,     5.7,     5.7,     5.7,
  4.98,    4.98,    4.98,    4.98,
  5.59,    5.59,    5.59,    5.59,
  5.32,    5.32,    5.32,    5.32,
  5.79,    5.79,    5.79,    5.79,
  5.63,    5.63,    5.63,    5.63,
  5.43,    5.43,    5.43,    5.43,
  5.68,    5.68,    5.68,    5.68,
  6.46,    6.46,    6.46,    6.46,
  6.39,    6.39,    6.39,    6.39,
  6.54,    6.54,    6.54,    6.54,
  6.43,    6.43,    6.43,    6.43,
  6.09,    6.09,    6.09,    6.09,
  5.96,    5.96,    5.96,    5.96,
  6.62,    6.62,    6.62,    6.62,
  6.36,    6.36,    6.36,    6.36,
  5.67,    5.67,    5.67,    5.67,
  5.61,    5.61,    5.61,    5.61,
  6.14,    6.14,    6.14,    6.14,
  5.91,    5.91,    5.91,    5.91,
  5.79,    5.79,    5.79,    5.79,
  6.27,    6.27,    6.27,    6.27,
  5.89,    5.89,    5.89,    5.89,
  6.08,    6.08,    6.08,    6.08,
  6.59,    6.59,    6.59,    6.59,
  7,       7,       7,       7,
  7.29,    7.29,    7.29,    7.29,
  7.75,    7.75,    7.75,    7.75,
  5.97,    5.97,    5.97,    5.97,
  6.62,    6.62,    6.62,    6.62,
  6.18,    6.18,    6.18,    6.18,
  6.01,    6.01,    6.01,    6.01,
  6.75,    6.75,    6.75,    6.75,
  6.26,    6.26,    6.26,    6.26,
  6.29,    6.29,    6.29,    6.29,
  6.64,    6.64,    6.64,    6.64,
  6.55,    6.55,    6.55,    6.55,
  6.11,    6.11,    6.11,    6.11,
  5.81,    5.81,    5.81,    5.81,
  6.31,    6.31,    6.31,    6.31,
  6.35,    6.35,    6.35,    6.35,
  6.25,    6.25,    6.25,    6.25,
  7.05,    7.05,    7.05,    7.05,
  6.95,    6.95,    6.95,    6.95,
  7.47,    7.47,    7.47,    7.47,
  7.27,    7.27,    7.27,    7.27,
  7.14,    7.14,    7.14,    7.14,
  7.15,    7.15,    7.15,    7.15,
  7.38,    7.38,    7.38,    7.38,
  6.96,    6.96,    6.96,    6.96,
  6.85,    6.85,    6.85,    6.85,
  7.11,    7.11,    7.11,    7.11,
  6.91,    6.91,    6.91,    6.91,
  6.31,    6.31,    6.31,    6.31,
  7.34,    7.34,    7.34,    7.34,
  6.85,    6.85,    6.85,    6.85,
  6.95,    6.95,    6.95,    6.95,
  7.19,    7.19,    7.19,    7.19,
  6.07,    6.07,    6.07,    6.07,
  6.1,     6.1,     6.1,     6.1,
  6.09,    6.09,    6.09,    6.09,
  5.27,    5.27,    5.27,    5.27,
  5.29,    5.29,    5.29,    5.29,
  5.68,    5.68,    5.68,    5.68,
  5.27,    5.27,    5.27,    5.27,
  5.82,    5.82,    5.82,    5.82,
  5.5,     5.5,     5.5,     5.5,
  5.82,    5.82,    5.82,    5.82,
  5.72,    5.72,    5.72,    5.72,
  5.87,    5.87,    5.87,    5.87,
  5.4,     5.4,     5.4,     5.4,
  5.83,    5.83,    5.83,    5.83,
  5.71,    5.71,    5.71,    5.71,
  4.87,    4.87,    4.87,    4.87,
  5.03,    5.03,    5.03,    5.03,
  5.45,    5.45,    5.45,    5.45,
  5.3,     5.3,     5.3,     5.3,
  5.13,    5.13,    5.13,    5.13,
  5.44,    5.44,    5.44,    5.44,
  4.47,    4.47,    4.47,    4.47,
  4.94,    4.94,    4.94,    4.94,
  4.84,    4.84,    4.84,    4.84,
  5.2,     5.2,     5.2,     5.2,
  5.11,    5.11,    5.11,    5.11,
  5.42,    5.42,    5.42,    5.42,
  4.75,    4.75,    4.75,    4.75,
  4.62,    4.62,    4.62,    4.62,
  4.9,     4.9,     4.9,     4.9,
  5.2,     5.2,     5.2,     5.2,
  4.64,    4.64,    4.64,    4.64,
  5,       5,       5,       5,
  4.68,    4.68,    4.68,    4.68,
  4.76,    4.76,    4.76,    4.76,
  4.09,    4.09,    4.09,    4.09,
  4.25,    4.25,    4.25,    4.25,
  4.36,    4.36,    4.36,    4.36,
  4.11,    4.11,    4.11,    4.11,
  4.25,    4.25,    4.25,    4.25,
  4.13,    4.13,    4.13,    4.13,
  4.59,    4.59,    4.59,    4.59,
  4.28,    4.28,    4.28,    4.28,
  3.68,    3.68,    3.68,    3.68,
  3.26,    3.26,    3.26,    3.26,
  4.75,    4.75,    4.75,    4.75,
  4.48,    4.48,    4.48,    4.48,
  4.65,    4.65,    4.65,    4.65,
  4.5,     4.5,     4.5,     4.5,
  4.29,    4.29,    4.29,    4.29,
  4.06,    4.06,    4.06,    4.06,
  3.67,    3.67,    3.67,    3.67,
  3.9,     3.9,     3.9,     3.9,
  4.2,     4.2,     4.2,     4.2,
  3.73,    3.73,    3.73,    3.73,
  3.36,    3.36,    3.36,    3.36,
  3.53,    3.53,    3.53,    3.53,
  3.52,    3.52,    3.52,    3.52,
  3.68,    3.68,    3.68,    3.68,
  3.93,    3.93,    3.93,    3.93,
  3.81,    3.81,    3.81,    3.81,
  3.54,    3.54,    3.54,    3.54,
  3.83,    3.83,    3.83,    3.83,
  3.77,    3.77,    3.77,    3.77,
  3.62,    3.62,    3.62,    3.62,
  3.77,    3.77,    3.77,    3.77,
  3.54,    3.54,    3.54,    3.54,
  3.46,    3.46,    3.46,    3.46,
  3.82,    3.82,    3.82,    3.82,
  3.27,    3.27,    3.27,    3.27,
  3.14,    3.14,    3.14,    3.14,
  3.41,    3.41,    3.41,    3.41,
  3.24,    3.24,    3.24,    3.24,
  2.94,    2.94,    2.94,    2.94,
  3.19,    3.19,    3.19,    3.19,
  2.76,    2.76,    2.76,    2.76,
  2.87,    2.87,    2.87,    2.87,
  2.97,    2.97,    2.97,    2.97,
  2.95,    2.95,    2.95,    2.95,
  2.93,    2.93,    2.93,    2.93,
  2.76,    2.76,    2.76,    2.76,
  3.08,    3.08,    3.08,    3.08,
  3.03,    3.03,    3.03,    3.03,
  2.96,    2.96,    2.96,    2.96,
  3.17,    3.17,    3.17,    3.17,
  3.12,    3.12,    3.12,    3.12,
  3.17,    3.17,    3.17,    3.17,
  2.91,    2.91,    2.91,    2.91,
  2.94,    2.94,    2.94,    2.94,
  3.54,    3.54,    3.54,    3.54,
  3.82,    3.82,    3.82,    3.82,
  3.54,    3.54,    3.54,    3.54,
  4.08,    4.08,    4.08,    4.08,
  3.98,    3.98,    3.98,    3.98,
  3.76,    3.76,    3.76,    3.76,
  3.61,    3.61,    3.61,    3.61,
  3.66,    3.66,    3.66,    3.66,
  3.73,    3.73,    3.73,    3.73,
  3.51,    3.51,    3.51,    3.51,
  3.66,    3.66,    3.66,    3.66,
  3.09,    3.09,    3.09,    3.09,
  3.4,     3.4,     3.4,     3.4,
  3.45,    3.45,    3.45,    3.45,
  3.82,    3.82,    3.82,    3.82,
  3.79,    3.79,    3.79,    3.79,
  4.03,    4.03,    4.03,    4.03,
  3.49,    3.49,    3.49,    3.49,
  4.2,     4.2,     4.2,     4.2,
  3.91,    3.91,    3.91,    3.91,
  3.84,    3.84,    3.84,    3.84,
  3.24,    3.24,    3.24,    3.24,
  2.51,    2.51,    2.51,    2.51,
  2.49,    2.49,    2.49,    2.49,
  2.62,    2.62,    2.62,    2.62,
  3.09,    3.09,    3.09,    3.09,
  2.66,    2.66,    2.66,    2.66,
  2.49,    2.49,    2.49,    2.49,
  2.59,    2.59,    2.59,    2.59,
  2.6,     2.6,     2.6,     2.6,
  2.45,    2.45,    2.45,    2.45,
  2.09,    2.09,    2.09,    2.09,
  2.32,    2.32,    2.32,    2.32,
  2.22,    2.22,    2.22,    2.22,
  2.03,    2.03,    2.03,    2.03,
  2.18,    2.18,    2.18,    2.18,
  1.83,    1.83,    1.83,    1.83,
  2.06,    2.06,    2.06,    2.06,
  2.21,    2.21,    2.21,    2.21,
  2.4,     2.4,     2.4,     2.4,
  2.32,    2.32,    2.32,    2.32,
  2.23,    2.23,    2.23,    2.23,
  2.22,    2.22,    2.22,    2.22,
  2.41,    2.41,    2.41,    2.41,
  2.52,    2.52,    2.52,    2.52,
  1.53,    1.53,    1.53,    1.53,
  1.44,    1.44,    1.44,    1.44,
  2.03,    2.03,    2.03,    2.03,
  2.36,    2.36,    2.36,    2.36,
  2.2,     2.2,     2.2,     2.2,
  2.44,    2.44,    2.44,    2.44,
  2.38,    2.38,    2.38,    2.38,
  2.32,    2.32,    2.32,    2.32,
  1.97,    1.97,    1.97,    1.97,
  1.83,    1.83,    1.83,    1.83,
  1.53,    1.53,    1.53,    1.53,
  1.31,    1.31,    1.31,    1.31,
  1.46,    1.46,    1.46,    1.46,
  1.37,    1.37,    1.37,    1.37,
  2.17,    2.17,    2.17,    2.17,
  1.57,    1.57,    1.57,    1.57,
  1.53,    1.53,    1.53,    1.53,
  1.86,    1.86,    1.86,    1.86,
  1.48,    1.48,    1.48,    1.48,
  1.53,    1.53,    1.53,    1.53,
  1.78,    1.78,    1.78,    1.78,
  2,       2,       2,       2,
  2.02,    2.02,    2.02,    2.02,
  1.83,    1.83,    1.83,    1.83,
  1.83,    1.83,    1.83,    1.83,
  1.76,    1.76,    1.76,    1.76,
  2.12,    2.12,    2.12,    2.12,
  2,       2,       2,       2,
  2.27,    2.27,    2.27,    2.27,
  2.12,    2.12,    2.12,    2.12,
  2.34,    2.34,    2.34,    2.34,
  2.63,    2.63,    2.63,    2.63,
  1.95,    1.95,    1.95,    1.95,
  1.69,    1.69,    1.69,    1.69,
  2.49,    2.49,    2.49,    2.49,
  2.25,    2.25,    2.25,    2.25,
  1.98,    1.98,    1.98,    1.98,
  1.66,    1.66,    1.66,    1.66,
  1.53,    1.53,    1.53,    1.53,
  1.95,    1.95,    1.95,    1.95,
  2.34,    2.34,    2.34,    2.34,
  2.5,     2.5,     2.5,     2.5,
  2.47,    2.47,    2.47,    2.47,
  2.5,     2.5,     2.5,     2.5,
  2.16,    2.16,    2.16,    2.16,
  2.16,    2.16,    2.16,    2.16,
  1.96,    1.96,    1.96,    1.96,
  2.01,    2.01,    2.01,    2.01,
  1.95,    1.95,    1.95,    1.95,
  1.89,    1.89,    1.89,    1.89,
  2.15,    2.15,    2.15,    2.15,
  2.25,    2.25,    2.25,    2.25,
  2.35,    2.35,    2.35,    2.35,
  2.47,    2.47,    2.47,    2.47,
  2.67,    2.67,    2.67,    2.67,
  3.13,    3.13,    3.13,    3.13,
  2.85,    2.85,    2.85,    2.85,
  2.69,    2.69,    2.69,    2.69,
  2.3,     2.3,     2.3,     2.3,
  2.31,    2.31,    2.31,    2.31,
  2.07,    2.07,    2.07,    2.07,
  2.51,    2.51,    2.51,    2.51,
  2.58,    2.58,    2.58,    2.58,
  2.14,    2.14,    2.14,    2.14,
  2.15,    2.15,    2.15,    2.15,
  2.08,    2.08,    2.08,    2.08,
  1.87,    1.87,    1.87,    1.87,
  1.78,    1.78,    1.78,    1.78,
  1.68,    1.68,    1.68,    1.68,
  2.12,    2.12,    2.12,    2.12,
  2.3,     2.3,     2.3,     2.3,
  1.95,    1.95,    1.95,    1.95,
  1.77,    1.77,    1.77,    1.77,
  1.98,    1.98,    1.98,    1.98,
  1.98,    1.98,    1.98,    1.98,
  2.03,    2.03,    2.03,    2.03,
  2.49,    2.49,    2.49,    2.49,
  2.57,    2.57,    2.57,    2.57,
  2.28,    2.28,    2.28,    2.28,
  1.78,    1.78,    1.78,    1.78,
  1.67,    1.67,    1.67,    1.67,
  2.35,    2.35,    2.35,    2.35,
  3.03,    3.03,    3.03,    3.03,
  2.23,    2.23,    2.23,    2.23,
  1.63,    1.63,    1.63,    1.63,
  1.36,    1.36,    1.36,    1.36,
  1.43,    1.43,    1.43,    1.43,
  1.43,    1.43,    1.43,    1.43,
  1.51,    1.51,    1.51,    1.51,
  1.73,    1.73,    1.73,    1.73,
  1.54,    1.54,    1.54,    1.54,
  1.55,    1.55,    1.55,    1.55,
  1.58,    1.58,    1.58,    1.58,
  1.72,    1.72,    1.72,    1.72,
  1.71,    1.71,    1.71,    1.71,
  1.36,    1.36,    1.36,    1.36,
  1.36,    1.36,    1.36,    1.36,
  1.66,    1.66,    1.66,    1.66,
  1.51,    1.51,    1.51,    1.51,
  1.49,    1.49,    1.49,    1.49,
  1,       1,       1,       1,
  0.85,    0.85,    0.85,    0.85,
  0.6,     0.6,     0.6,     0.6,
  1.04,    1.04,    1.04,    1.04,
  1.21,    1.21,    1.21,    1.21,
  1.74,    1.74,    1.74,    1.74,
  0.81,    0.81,    0.81,    0.81,
  0.76,    0.76,    0.76,    0.76,
  0.8,     0.8,     0.8,     0.8,
  0.82,    0.82,    0.82,    0.82,
  1.14,    1.14,    1.14,    1.14,
  0.97,    0.97,    0.97,    0.97,
  1.19,    1.19,    1.19,    1.19,
  0.89,    0.89,    0.89,    0.89,
  0.98,    0.98,    0.98,    0.98,
  0.98,    0.98,    0.98,    0.98,
  0.77,    0.77,    0.77,    0.77,
  0.74,    0.74,    0.74,    0.74,
  1.26,    1.26,    1.26,    1.26,
  1.23,    1.23,    1.23,    1.23,
  1.13,    1.13,    1.13,    1.13,
  0.88,    0.88,    0.88,    0.88,
  0.57,    0.57,    0.57,    0.57,
  0.81,    0.81,    0.81,    0.81,
  0.83,    0.83,    0.83,    0.83,
  0.68,    0.68,    0.68,    0.68,
  0.78,    0.78,    0.78,    0.78,
  0.77,    0.77,    0.77,    0.77,
  0.58,    0.58,    0.58,    0.58,
  0.75,    0.75,    0.75,    0.75,
  0.44,    0.44,    0.44,    0.44,
  0.41,    0.41,    0.41,    0.41,
  0.59,    0.59,    0.59,    0.59,
  1.12,    1.12,    1.12,    1.12,
  1.13,    1.13,    1.13,    1.13,
  0.88,    0.88,    0.88,    0.88,
  0.91,    0.91,    0.91,    0.91,
  1.03,    1.03,    1.03,    1.03,
  1.09,    1.09,    1.09,    1.09,
  0.98,    0.98,    0.98,    0.98,
  0.93,    0.93,    0.93,    0.93,
  0.86,    0.86,    0.86,    0.86,
  0.75,    0.75,    0.75,    0.75,
  1.12,    1.12,    1.12,    1.12,
  1.26,    1.26,    1.26,    1.26,
  1.38,    1.38,    1.38,    1.38,
  0.92,    0.92,    0.92,    0.92,
  1.18,    1.18,    1.18,    1.18,
  1.28,    1.28,    1.28,    1.28,
  1.46,    1.46,    1.46,    1.46,
  1.37,    1.37,    1.37,    1.37,
  1.15,    1.15,    1.15,    1.15,
  1.46,    1.46,    1.46,    1.46,
  1.51,    1.51,    1.51,    1.51,
  1.51,    1.51,    1.51,    1.51,
  1.42,    1.42,    1.42,    1.42,
  1.72,    1.72,    1.72,    1.72,
  1.52,    1.52,    1.52,    1.52,
  2.02,    2.02,    2.02,    2.02,
  1.83,    1.83,    1.83,    1.83,
  1.76,    1.76,    1.76,    1.76,
  1.6,     1.6,     1.6,     1.6,
  1.88,    1.88,    1.88,    1.88,
  2.07,    2.07,    2.07,    2.07,
  2.17,    2.17,    2.17,    2.17,
  2.17,    2.17,    2.17,    2.17,
  2.27,    2.27,    2.27,    2.27,
  2.65,    2.65,    2.65,    2.65,
  2.67,    2.67,    2.67,    2.67,
  2.12,    2.12,    2.12,    2.12,
  2.26,    2.26,    2.26,    2.26,
  2.11,    2.11,    2.11,    2.11,
  2.23,    2.23,    2.23,    2.23,
  2.88,    2.88,    2.88,    2.88,
  3.22,    3.22,    3.22,    3.22,
  2.89,    2.89,    2.89,    2.89,
  2.65,    2.65,    2.65,    2.65,
  2.71,    2.71,    2.71,    2.71,
  2.94,    2.94,    2.94,    2.94,
  3.08,    3.08,    3.08,    3.08,
  3.09,    3.09,    3.09,    3.09,
  2.62,    2.62,    2.62,    2.62,
  3.06,    3.06,    3.06,    3.06,
  3.4,     3.4,     3.4,     3.4,
  3.48,    3.48,    3.48,    3.48,
  3.41,    3.41,    3.41,    3.41,
  3.62,    3.62,    3.62,    3.62,
  4.18,    4.18,    4.18,    4.18,
  3.46,    3.46,    3.46,    3.46,
  3.51,    3.51,    3.51,    3.51,
  3.6,     3.6,     3.6,     3.6,
  3.58,    3.58,    3.58,    3.58,
  3.85,    3.85,    3.85,    3.85,
  3.33,    3.33,    3.33,    3.33,
  3.27,    3.27,    3.27,    3.27,
  3.36,    3.36,    3.36,    3.36,
  3.31,    3.31,    3.31,    3.31,
  3.51,    3.51,    3.51,    3.51,
  3.07,    3.07,    3.07,    3.07,
  3.21,    3.21,    3.21,    3.21,
  2.99,    2.99,    2.99,    2.99,
  3.19,    3.19,    3.19,    3.19,
  3.09,    3.09,    3.09,    3.09,
  2.77,    2.77,    2.77,    2.77,
  2.55,    2.55,    2.55,    2.55,
  2.94,    2.94,    2.94,    2.94,
  2.63,    2.63,    2.63,    2.63,
  3.2,     3.2,     3.2,     3.2,
  3.39,    3.39,    3.39,    3.39,
  2.92,    2.92,    2.92,    2.92,
  3.54,    3.54,    3.54,    3.54,
  3.68,    3.68,    3.68,    3.68,
  4.02,    4.02,    4.02,    4.02,
  3.78,    3.78,    3.78,    3.78,
  4.09,    4.09,    4.09,    4.09,
  4.23,    4.23,    4.23,    4.23,
  5.32,    5.32,    5.32,    5.32,
  5.38,    5.38,    5.38,    5.38,
  5.91,    5.91,    5.91,    5.91,
  5.64,    5.64,    5.64,    5.64,
  5.38,    5.38,    5.38,    5.38,
  5.69,    5.69,    5.69,    5.69,
  5.07,    5.07,    5.07,    5.07,
  5.77,    5.77,    5.77,    5.77,
  5.42,    5.42,    5.42,    5.42,
  6.66,    6.66,    6.66,    6.66,
  7.02,    7.02,    7.02,    7.02,
  5.38,    5.38,    5.38,    5.38,
  6.2,     6.2,     6.2,     6.2,
  6.8,     6.8,     6.8,     6.8,
  6,       6,       6,       6,
  5.89,    5.89,    5.89,    5.89,
  6.46,    6.46,    6.46,    6.46,
  5.75,    5.75,    5.75,    5.75,
  5.16,    5.16,    5.16,    5.16,
  5.17,    5.17,    5.17,    5.17,
  5.08,    5.08,    5.08,    5.08,
  4.79,    4.79,    4.79,    4.79,
  4.92,    4.92,    4.92,    4.92,
  4.6,     4.6,     4.6,     4.6,
  4.79,    4.79,    4.79,    4.79,
  4.56,    4.56,    4.56,    4.56,
  4.8,     4.8,     4.8,     4.8,
  4.69,    4.69,    4.69,    4.69,
  4.55,    4.55,    4.55,    4.55,
  4.84,    4.84,    4.84,    4.84,
  4.53,    4.53,    4.53,    4.53,
  4.45,    4.45,    4.45,    4.45,
  5.01,    5.01,    5.01,    5.01,
  4.67,    4.67,    4.67,    4.67,
  4.73,    4.73,    4.73,    4.73,
  4.28,    4.28,    4.28,    4.28,
  4.16,    4.16,    4.16,    4.16,
  3.87,    3.87,    3.87,    3.87,
  3.33,    3.33,    3.33,    3.33,
  4.64,    4.64,    4.64,    4.64,
  4.8,     4.8,     4.8,     4.8,
  6.84,    6.84,    6.84,    6.84,
  5.55,    5.55,    5.55,    5.55,
  5.74,    5.74,    5.74,    5.74,
  5.43,    5.43,    5.43,    5.43,
  6.61,    6.61,    6.61,    6.61,
  7.1,     7.1,     7.1,     7.1,
  6.3,     6.3,     6.3,     6.3,
  6.49,    6.49,    6.49,    6.49,
  6.7,     6.7,     6.7,     6.7,
  6.77,    6.77,    6.77,    6.77,
  6.88,    6.88,    6.88,    6.88,
  6.02,    6.02,    6.02,    6.02,
  6.27,    6.27,    6.27,    6.27,
  6.66,    6.66,    6.66,    6.66,
  6.87,    6.87,    6.87,    6.87,
  7.19,    7.19,    7.19,    7.19,
  6.36,    6.36,    6.36,    6.36,
  6.71,    6.71,    6.71,    6.71,
  7.04,    7.04,    7.04,    7.04,
  6.74,    6.74,    6.74,    6.74,
  7.34,    7.34,    7.34,    7.34,
  6.85,    6.85,    6.85,    6.85,
  6.91,    6.91,    6.91,    6.91,
  7.41,    7.41,    7.41,    7.41,
  6.86,    6.86,    6.86,    6.86,
  6.64,    6.64,    6.64,    6.64,
  6.97,    6.97,    6.97,    6.97,
  7.6,     7.6,     7.6,     7.6,
  7.15,    7.15,    7.15,    7.15,
  6.57,    6.57,    6.57,    6.57,
  6.74,    6.74,    6.74,    6.74,
  6.77,    6.77,    6.77,    6.77,
  7.53,    7.53,    7.53,    7.53,
  7.13,    7.13,    7.13,    7.13,
  6.44,    6.44,    6.44,    6.44,
  6.66,    6.66,    6.66,    6.66,
  6.54,    6.54,    6.54,    6.54,
  6.01,    6.01,    6.01,    6.01,
  6.09,    6.09,    6.09,    6.09,
  5.93,    5.93,    5.93,    5.93,
  6.33,    6.33,    6.33,    6.33,
  5.86,    5.86,    5.86,    5.86,
  6.14,    6.14,    6.14,    6.14,
  6.24,    6.24,    6.24,    6.24,
  4.74,    4.74,    4.74,    4.74,
  5.02,    5.02,    5.02,    5.02,
  4.55,    4.55,    4.55,    4.55,
  4.56,    4.56,    4.56,    4.56,
  4.24,    4.24,    4.24,    4.24,
  3.86,    3.86,    3.86,    3.86,
  3.84,    3.84,    3.84,    3.84,
  3.67,    3.67,    3.67,    3.67,
  3.27,    3.27,    3.27,    3.27,
  3.06,    3.06,    3.06,    3.06,
  2.95,    2.95,    2.95,    2.95,
  2.31,    2.31,    2.31,    2.31,
  2.56,    2.56,    2.56,    2.56,
  2.17,    2.17,    2.17,    2.17,
  2.44,    2.44,    2.44,    2.44,
  2.89,    2.89,    2.89,    2.89,
  3.85,    3.85,    3.85,    3.85,
  3.53,    3.53,    3.53,    3.53,
  1.95,    1.95,    1.95,    1.95,
  1.83,    1.83,    1.83,    1.83,
  2.44,    2.44,    2.44,    2.44,
  2.47,    2.47,    2.47,    2.47,
  2.26,    2.26,    2.26,    2.26,
  2.42,    2.42,    2.42,    2.42,
  2.5,     2.5,     2.5,     2.5,
  2.58,    2.58,    2.58,    2.58,
  2.55,    2.55,    2.55,    2.55,
  2.76,    2.76,    2.76,    2.76,
  2.72,    2.72,    2.72,    2.72,
  2.72,    2.72,    2.72,    2.72,
  2.76,    2.76,    2.76,    2.76,
  3.02,    3.02,    3.02,    3.02,
  2.64,    2.64,    2.64,    2.64,
  2.05,    2.05,    2.05,    2.05,
  2.17,    2.17,    2.17,    2.17,
  2.58,    2.58,    2.58,    2.58,
  2.17,    2.17,    2.17,    2.17,
  2.17,    2.17,    2.17,    2.17,
  2.17,    2.17,    2.17,    2.17,
  2.13,    2.13,    2.13,    2.13,
  1.91,    1.91,    1.91,    1.91,
  2.32,    2.32,    2.32,    2.32,
  2.3,     2.3,     2.3,     2.3,
  2.42,    2.42,    2.42,    2.42,
  2.19,    2.19,    2.19,    2.19,
  2.43,    2.43,    2.43,    2.43,
  2,       2,       2,       2,
  2,       2,       2,       2,
  2.17,    2.17,    2.17,    2.17,
  2.77,    2.77,    2.77,    2.77,
  2.56,    2.56,    2.56,    2.56,
  2.25,    2.25,    2.25,    2.25,
  2.4,     2.4,     2.4,     2.4,
  1.97,    1.97,    1.97,    1.97,
  1.72,    1.72,    1.72,    1.72,
  1.49,    1.49,    1.49,    1.49,
  1.95,    1.95,    1.95,    1.95,
  1.78,    1.78,    1.78,    1.78,
  1.85,    1.85,    1.85,    1.85,
  1.95,    1.95,    1.95,    1.95,
  1.98,    1.98,    1.98,    1.98,
  2.23,    2.23,    2.23,    2.23,
  2.24,    2.24,    2.24,    2.24,
  2.06,    2.06,    2.06,    2.06,
  2.38,    2.38,    2.38,    2.38,
  2.14,    2.14,    2.14,    2.14,
  1.63,    1.63,    1.63,    1.63,
  1.52,    1.52,    1.52,    1.52,
  1.53,    1.53,    1.53,    1.53,
  1.67,    1.67,    1.67,    1.67,
  1.8,     1.8,     1.8,     1.8,
  1.86,    1.86,    1.86,    1.86,
  1.91,    1.91,    1.91,    1.91,
  2.19,    2.19,    2.19,    2.19,
  1.45,    1.45,    1.45,    1.45,
  1.73,    1.73,    1.73,    1.73,
  1.74,    1.74,    1.74,    1.74,
  1.96,    1.96,    1.96,    1.96,
  1.95,    1.95,    1.95,    1.95,
  1.99,    1.99,    1.99,    1.99,
  2.21,    2.21,    2.21,    2.21,
  2.22,    2.22,    2.22,    2.22,
  2,       2,       2,       2,
  2.14,    2.14,    2.14,    2.14,
  2.37,    2.37,    2.37,    2.37,
  2.06,    2.06,    2.06,    2.06,
  2.26,    2.26,    2.26,    2.26,
  1.76,    1.76,    1.76,    1.76,
  2.18,    2.18,    2.18,    2.18,
  2.17,    2.17,    2.17,    2.17,
  2.3,     2.3,     2.3,     2.3,
  2.03,    2.03,    2.03,    2.03,
  2.22,    2.22,    2.22,    2.22,
  2.21,    2.21,    2.21,    2.21,
  3.18,    3.18,    3.18,    3.18,
  3.08,    3.08,    3.08,    3.08,
  3.41,    3.41,    3.41,    3.41,
  3.35,    3.35,    3.35,    3.35,
  2.84,    2.84,    2.84,    2.84,
  2.43,    2.43,    2.43,    2.43,
  3.04,    3.04,    3.04,    3.04,
  2.78,    2.78,    2.78,    2.78,
  2.85,    2.85,    2.85,    2.85,
  3.32,    3.32,    3.32,    3.32,
  3.44,    3.44,    3.44,    3.44,
  3.8,     3.8,     3.8,     3.8,
  4.08,    4.08,    4.08,    4.08,
  3.97,    3.97,    3.97,    3.97,
  4.59,    4.59,    4.59,    4.59,
  4.18,    4.18,    4.18,    4.18,
  5.11,    5.11,    5.11,    5.11,
  4.95,    4.95,    4.95,    4.95,
  4.86,    4.86,    4.86,    4.86,
  4.67,    4.67,    4.67,    4.67,
  4.37,    4.37,    4.37,    4.37,
  3.8,     3.8,     3.8,     3.8,
  3.55,    3.55,    3.55,    3.55,
  3.36,    3.36,    3.36,    3.36,
  3.13,    3.13,    3.13,    3.13,
  3.5,     3.5,     3.5,     3.5,
  3.47,    3.47,    3.47,    3.47,
  2.91,    2.91,    2.91,    2.91,
  2.81,    2.81,    2.81,    2.81,
  2.79,    2.79,    2.79,    2.79,
  2.35,    2.35,    2.35,    2.35,
  2.25,    2.25,    2.25,    2.25,
  2.25,    2.25,    2.25,    2.25,
  2.77,    2.77,    2.77,    2.77,
  3.1,     3.1,     3.1,     3.1,
  2.29,    2.29,    2.29,    2.29,
  2.07,    2.07,    2.07,    2.07,
  2.21,    2.21,    2.21,    2.21,
  2.46,    2.46,    2.46,    2.46,
  2.29,    2.29,    2.29,    2.29,
  2.25,    2.25,    2.25,    2.25,
  2.44,    2.44,    2.44,    2.44,
  2.12,    2.12,    2.12,    2.12,
  2.1,     2.1,     2.1,     2.1,
  2.16,    2.16,    2.16,    2.16,
  2.26,    2.26,    2.26,    2.26,
  1.77,    1.77,    1.77,    1.77,
  1.79,    1.79,    1.79,    1.79,
  2.17,    2.17,    2.17,    2.17,
  2.5,     2.5,     2.5,     2.5,
  2.3,     2.3,     2.3,     2.3,
  2.13,    2.13,    2.13,    2.13,
  1.82,    1.82,    1.82,    1.82,
  2.54,    2.54,    2.54,    2.54,
  2.52,    2.52,    2.52,    2.52,
  1.92,    1.92,    1.92,    1.92,
  1.66,    1.66,    1.66,    1.66,
  1.95,    1.95,    1.95,    1.95,
  2.26,    2.26,    2.26,    2.26,
  2.32,    2.32,    2.32,    2.32,
  2.63,    2.63,    2.63,    2.63,
  2.38,    2.38,    2.38,    2.38,
  2.53,    2.53,    2.53,    2.53,
  2.55,    2.55,    2.55,    2.55,
  2.5,     2.5,     2.5,     2.5,
  2.76,    2.76,    2.76,    2.76,
  2.59,    2.59,    2.59,    2.59,
  2.54,    2.54,    2.54,    2.54,
  2.69,    2.69,    2.69,    2.69,
  2.57,    2.57,    2.57,    2.57,
  2.62,    2.62,    2.62,    2.62,
  2.58,    2.58,    2.58,    2.58,
  2.32,    2.32,    2.32,    2.32,
  2.54,    2.54,    2.54,    2.54,
  2.23,    2.23,    2.23,    2.23,
  2.74,    2.74,    2.74,    2.74,
  2.36,    2.36,    2.36,    2.36,
  3.28,    3.28,    3.28,    3.28,
  2.88,    2.88,    2.88,    2.88,
  2.55,    2.55,    2.55,    2.55,
  2.61,    2.61,    2.61,    2.61,
  1.74,    1.74,    1.74,    1.74,
  1.94,    1.94,    1.94,    1.94,
  1.61,    1.61,    1.61,    1.61,
  1.89,    1.89,    1.89,    1.89,
  2.16,    2.16,    2.16,    2.16,
  1.97,    1.97,    1.97,    1.97,
  2.44,    2.44,    2.44,    2.44,
  2.47,    2.47,    2.47,    2.47,
  2.67,    2.67,    2.67,    2.67,
  2.67,    2.67,    2.67,    2.67,
  2.53,    2.53,    2.53,    2.53,
  2.64,    2.64,    2.64,    2.64,
  3.09,    3.09,    3.09,    3.09,
  3.09,    3.09,    3.09,    3.09,
  3.12,    3.12,    3.12,    3.12,
  3.3,     3.3,     3.3,     3.3,
  3.1,     3.1,     3.1,     3.1,
  3.22,    3.22,    3.22,    3.22,
  3.27,    3.27,    3.27,    3.27,
  3.47,    3.47,    3.47,    3.47,
  3.21,    3.21,    3.21,    3.21,
  3.04,    3.04,    3.04,    3.04,
  3.07,    3.07,    3.07,    3.07,
  3.39,    3.39,    3.39,    3.39,
  2.99,    2.99,    2.99,    2.99,
  3.15,    3.15,    3.15,    3.15,
  3.26,    3.26,    3.26,    3.26,
  3.03,    3.03,    3.03,    3.03,
  3.48,    3.48,    3.48,    3.48,
  3.29,    3.29,    3.29,    3.29,
  3.9,     3.9,     3.9,     3.9,
  3.76,    3.76,    3.76,    3.76,
  3.64,    3.64,    3.64,    3.64,
  3.57,    3.57,    3.57,    3.57,
  3.3,     3.3,     3.3,     3.3,
  3.87,    3.87,    3.87,    3.87,
  3.72,    3.72,    3.72,    3.72,
  3.31,    3.31,    3.31,    3.31,
  3.36,    3.36,    3.36,    3.36,
  3.77,    3.77,    3.77,    3.77,
  3.75,    3.75,    3.75,    3.75,
  3.48,    3.48,    3.48,    3.48,
  4.08,    4.08,    4.08,    4.08,
  4.09,    4.09,    4.09,    4.09,
  4.1,     4.1,     4.1,     4.1,
  3.84,    3.84,    3.84,    3.84,
  4.2,     4.2,     4.2,     4.2,
  4.71,    4.71,    4.71,    4.71,
  4.53,    4.53,    4.53,    4.53,
  4.09,    4.09,    4.09,    4.09,
  4.53,    4.53,    4.53,    4.53,
  4.32,    4.32,    4.32,    4.32,
  4.17,    4.17,    4.17,    4.17,
  3.89,    3.89,    3.89,    3.89,
  4.25,    4.25,    4.25,    4.25,
  4.71,    4.71,    4.71,    4.71,
  4.52,    4.52,    4.52,    4.52,
  4.46,    4.46,    4.46,    4.46,
  4.47,    4.47,    4.47,    4.47,
  4.29,    4.29,    4.29,    4.29,
  4.8,     4.8,     4.8,     4.8,
  4.5,     4.5,     4.5,     4.5,
  4.94,    4.94,    4.94,    4.94,
  4.21,    4.21,    4.21,    4.21,
  4.05,    4.05,    4.05,    4.05,
  3.94,    3.94,    3.94,    3.94,
  3.75,    3.75,    3.75,    3.75,
  3.25,    3.25,    3.25,    3.25,
  3.41,    3.41,    3.41,    3.41,
  2.81,    2.81,    2.81,    2.81,
  2.55,    2.55,    2.55,    2.55,
  2.07,    2.07,    2.07,    2.07,
  1.82,    1.82,    1.82,    1.82,
  2.01,    2.01,    2.01,    2.01,
  1.72,    1.72,    1.72,    1.72,
  1.72,    1.72,    1.72,    1.72,
  1.5,     1.5,     1.5,     1.5,
  1.57,    1.57,    1.57,    1.57,
  1.72,    1.72,    1.72,    1.72,
  1.69,    1.69,    1.69,    1.69,
  1.68,    1.68,    1.68,    1.68,
  1.39,    1.39,    1.39,    1.39,
  1.66,    1.66,    1.66,    1.66,
  1.62,    1.62,    1.62,    1.62,
  1.83,    1.83,    1.83,    1.83,
  1.79,  1.79,  1.79,   1.79 ;

 PSurf =
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  104200,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103900,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103200,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  103500,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  100200,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99600,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99500,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  103000,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  102500,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100300,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101700,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102400,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103800,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103400,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  103100,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102600,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  102200,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  101000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  100000,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  98900,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99300,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99100,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99400,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  99700,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101200,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  102000,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102100,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  102300,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101900,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  101500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  100100,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102800,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  102900,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  103300,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  102700,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  101300,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  99900,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101100,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101600,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101800,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  101400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  100400,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  99800,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100600,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100800,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100900,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100700,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500,
  100500 ;

 LWdown =
  187.8,
  186.9,
  186.7,
  187.3,
  187.3,
  187.5,
  187.2,
  187,
  186.4,
  186.3,
  186.3,
  186.3,
  186.6,
  187.2,
  186.9,
  187.4,
  187.6,
  187.8,
  186.8,
  185.8,
  186.4,
  188,
  188.3,
  189.1,
  185.8,
  178.2,
  189.7,
  192.7,
  192.2,
  191.6,
  191.8,
  248,
  208.4,
  193.5,
  192.5,
  192.3,
  192,
  192.1,
  192,
  191.3,
  191.3,
  193.2,
  191.7,
  191.5,
  191.1,
  191,
  192,
  191.9,
  190.7,
  191.6,
  192.2,
  194.1,
  192.5,
  193.5,
  193,
  193.6,
  194.1,
  195.1,
  193.9,
  194.7,
  196,
  193.3,
  191.7,
  192,
  191.6,
  191.5,
  189.5,
  188.3,
  187.8,
  188.7,
  187.7,
  189,
  189.4,
  186.5,
  197.3,
  199.3,
  198.5,
  196.7,
  196.5,
  249.2,
  211.6,
  195.5,
  195.3,
  194.7,
  194.5,
  194.3,
  193.7,
  193.6,
  192.9,
  192.8,
  192.4,
  192.1,
  192.3,
  192,
  192.2,
  192.7,
  194,
  194.5,
  196,
  197.6,
  197.6,
  197.3,
  198.2,
  203.5,
  218.6,
  234.4,
  233.9,
  232.7,
  238.8,
  247.9,
  249.8,
  253.9,
  247.9,
  253.6,
  256.7,
  260,
  256.8,
  258.1,
  259.1,
  263.5,
  265.5,
  270,
  269.3,
  258,
  243.6,
  241.8,
  285,
  306.9,
  290.2,
  262,
  255,
  268.7,
  257.8,
  257.3,
  267.1,
  288.2,
  284.3,
  285.3,
  277.9,
  278.4,
  281.4,
  282.3,
  282.8,
  283.3,
  283.8,
  284.1,
  284.3,
  284.6,
  285.4,
  285.8,
  285.9,
  286.2,
  286.4,
  286.6,
  286.4,
  286.2,
  286.2,
  285,
  285.1,
  284.6,
  284.3,
  284.9,
  283.9,
  284,
  284.2,
  283.6,
  283.9,
  285.5,
  287.1,
  289.3,
  289.4,
  293.3,
  295.3,
  297.1,
  297.1,
  308.1,
  298.5,
  294.4,
  291.5,
  291.4,
  294.7,
  299.4,
  298.8,
  298.9,
  298.4,
  297.9,
  297.9,
  296.4,
  296.1,
  293.2,
  263.2,
  286,
  273.2,
  282.9,
  296.7,
  297.2,
  297.4,
  296.9,
  296.2,
  295.8,
  291.8,
  260.6,
  244.4,
  268.5,
  289,
  289.7,
  287.5,
  287.9,
  288,
  287.2,
  284.3,
  279.1,
  286.7,
  287.9,
  290.1,
  292.4,
  292.2,
  291.1,
  285.1,
  249.8,
  208.7,
  205.1,
  205.3,
  268.1,
  229,
  210.1,
  210.1,
  211.6,
  212.4,
  210.5,
  208.5,
  207.5,
  206.7,
  207.4,
  205,
  202.8,
  201.7,
  237.1,
  240.6,
  233.8,
  223.6,
  205.7,
  211.2,
  270.1,
  272.5,
  270.2,
  274.2,
  276,
  279.2,
  280.1,
  275.7,
  277.4,
  272.9,
  271.8,
  277.7,
  277.9,
  278.6,
  279.3,
  278.7,
  275.8,
  274.6,
  270.7,
  268.7,
  264.2,
  246.6,
  207.9,
  208.1,
  210.9,
  207.7,
  205.6,
  203.2,
  286.4,
  233.3,
  204.1,
  203.3,
  203.9,
  204,
  204.1,
  203.5,
  203.4,
  215.8,
  246.2,
  268.8,
  269.2,
  273.5,
  279.1,
  271.9,
  278.5,
  275.3,
  280.9,
  280.4,
  280.3,
  281.4,
  283.1,
  283.6,
  284.2,
  281.9,
  281.7,
  283.3,
  284.5,
  284.8,
  286.2,
  287.1,
  287.1,
  286.1,
  285.5,
  285.1,
  285.4,
  285.6,
  285.9,
  271.6,
  280.3,
  282.2,
  282.1,
  269.3,
  270.5,
  260.3,
  245.2,
  217.7,
  265.4,
  235.9,
  221.2,
  222.8,
  223.3,
  223.4,
  221.3,
  218.1,
  217.9,
  217,
  235.9,
  266.6,
  270.4,
  253.9,
  241.8,
  240.9,
  241.3,
  254.4,
  245.9,
  257.1,
  252.2,
  256.7,
  256.8,
  248.2,
  237.2,
  233.5,
  224.5,
  216.5,
  215,
  214.7,
  215.3,
  227.5,
  243.2,
  250.7,
  256.6,
  264.5,
  265.5,
  268,
  270.7,
  272.4,
  272.6,
  272,
  263.5,
  252.2,
  259.3,
  268.2,
  256.1,
  247.1,
  248.2,
  251.1,
  232.9,
  228.7,
  226.1,
  221.5,
  220.5,
  220.5,
  221.4,
  223.2,
  223.3,
  228.7,
  237.3,
  241.5,
  241.7,
  247.1,
  246.7,
  241.3,
  234.5,
  232.3,
  238.4,
  240.4,
  241.3,
  240.6,
  246.4,
  244.9,
  241.1,
  243.4,
  232.8,
  225.8,
  231.7,
  249.8,
  260.3,
  265.2,
  269.6,
  269.9,
  269.7,
  265.9,
  261.9,
  254.8,
  247.3,
  250,
  250.1,
  248.9,
  253.4,
  245.3,
  239.7,
  240.3,
  264.2,
  250.3,
  235.8,
  253.2,
  269.6,
  276.1,
  281.7,
  283.8,
  285.3,
  285.8,
  286.1,
  287.2,
  288.2,
  289.5,
  290.1,
  289.8,
  289.6,
  289.8,
  290.5,
  290.9,
  291.5,
  291.7,
  292.2,
  292.4,
  292.5,
  292.1,
  291.5,
  290.6,
  289.2,
  288.8,
  288.3,
  287.8,
  287.9,
  288,
  287.4,
  286.9,
  287.6,
  287.5,
  287.1,
  286.6,
  287.6,
  282,
  281.1,
  278.8,
  284.9,
  285.7,
  287.8,
  289,
  298.2,
  292.8,
  289.8,
  290.1,
  289.7,
  290.2,
  290.6,
  291,
  290.9,
  290.7,
  291.6,
  290.9,
  291.2,
  290.8,
  291.4,
  291.5,
  291.5,
  291.1,
  291.3,
  291.5,
  291,
  290.6,
  290.3,
  289.6,
  289,
  288.2,
  287.9,
  288,
  288.1,
  287.7,
  288,
  288.2,
  288,
  288.4,
  288.1,
  288.4,
  288.8,
  289.1,
  289.8,
  290.1,
  290.4,
  290.2,
  289.8,
  288.8,
  288.2,
  285.6,
  285.2,
  284.3,
  299,
  279.6,
  281,
  285.5,
  285.1,
  284.7,
  283.4,
  270.1,
  229.2,
  230.7,
  231.8,
  233.1,
  233.8,
  233.7,
  233.8,
  234,
  233.8,
  233.8,
  234.2,
  234.3,
  235.3,
  236.3,
  246.5,
  259,
  286,
  296.6,
  298.5,
  303.7,
  300.6,
  302.5,
  304.8,
  313.5,
  311.1,
  311.8,
  312.9,
  312.1,
  315.3,
  317.5,
  317.8,
  318.5,
  320,
  318.3,
  316.6,
  318,
  320.6,
  319,
  319,
  320.2,
  342.5,
  329.7,
  323.7,
  321.3,
  321.9,
  323.2,
  323.2,
  323.3,
  324.2,
  325.2,
  325.3,
  325.8,
  325.3,
  325.3,
  325.2,
  325.2,
  325.3,
  325.8,
  325.8,
  326,
  325.9,
  326.2,
  326.7,
  326.2,
  325.9,
  325.8,
  325.8,
  326.1,
  326.1,
  325.7,
  325.1,
  325.5,
  325.3,
  325,
  325,
  325.5,
  324.2,
  325.6,
  312.5,
  269.1,
  262.4,
  264.3,
  261.8,
  269.3,
  270.9,
  271.1,
  271.3,
  271.4,
  352.7,
  307.6,
  277.7,
  272.5,
  273,
  275.7,
  275.1,
  276.6,
  276,
  278.3,
  277.7,
  277.9,
  277.9,
  274.2,
  267.3,
  263.7,
  262.4,
  264.2,
  264.3,
  264.3,
  263.3,
  262.5,
  262.5,
  259.9,
  259.1,
  258.9,
  257.9,
  257.9,
  258.2,
  259.3,
  260.1,
  258.3,
  258.3,
  258.3,
  258.8,
  257.9,
  260.5,
  265.2,
  268.5,
  273.4,
  275.8,
  274.1,
  270.4,
  278.5,
  282.2,
  281.6,
  282,
  278.9,
  275.5,
  327.4,
  283.8,
  266.6,
  261.8,
  260.5,
  259.4,
  260.8,
  258.4,
  253.5,
  251.3,
  249.6,
  246.3,
  245.4,
  246.3,
  244.8,
  241.3,
  241.7,
  242.2,
  241.5,
  241,
  240.2,
  238.6,
  236.6,
  235,
  235.1,
  234.6,
  234,
  234.2,
  233.3,
  233.6,
  232.8,
  231.7,
  231.8,
  232.1,
  231.6,
  230.6,
  230.9,
  233.2,
  235.8,
  237.5,
  237.8,
  229.7,
  240.4,
  245.1,
  247.4,
  247.2,
  248.8,
  250.1,
  288.4,
  259.3,
  252.5,
  254.4,
  251.5,
  249.3,
  248.3,
  248.2,
  246.9,
  245.2,
  245.8,
  244.7,
  245.1,
  245.3,
  245.3,
  246.3,
  246.9,
  245.6,
  244.4,
  241.7,
  241.3,
  241.9,
  243.3,
  242.5,
  240.9,
  239.4,
  238.8,
  238.7,
  239.3,
  239.1,
  239.1,
  238.3,
  238,
  238,
  236.7,
  236,
  237.3,
  240.6,
  243.6,
  246.4,
  248.3,
  240.6,
  253.9,
  257.1,
  258.1,
  260.5,
  258.9,
  260.6,
  303.3,
  263.9,
  250.4,
  249.6,
  248.4,
  247.8,
  246,
  246,
  245.4,
  244.6,
  244.7,
  245,
  246.9,
  247.3,
  245.8,
  245.1,
  245,
  244.2,
  245.2,
  243.8,
  244.3,
  244.7,
  243.5,
  244.4,
  242.9,
  245.2,
  245.2,
  245.5,
  246.3,
  246.6,
  246.3,
  246.6,
  248.2,
  249.5,
  249.2,
  247.2,
  248.7,
  252,
  255.2,
  257.5,
  259.3,
  250.9,
  261.2,
  265.5,
  265,
  264.4,
  263.6,
  263.4,
  282.5,
  267.1,
  264,
  263.4,
  264,
  265.5,
  267.2,
  268.9,
  270.3,
  297.8,
  334,
  339.4,
  343.8,
  344.9,
  342.8,
  342,
  341.8,
  340.8,
  341.2,
  340.2,
  338.5,
  340.3,
  340.6,
  339.5,
  338.9,
  339.2,
  339.3,
  339.4,
  339.3,
  339.3,
  340.3,
  340.5,
  340.9,
  341.8,
  342.3,
  342.4,
  342.3,
  342.6,
  342.4,
  341.8,
  341.3,
  341.7,
  343,
  343.2,
  344.3,
  343.8,
  343.6,
  342.5,
  347.5,
  343.3,
  340.7,
  340,
  339.9,
  339.4,
  339.5,
  338.8,
  338.4,
  337.9,
  337.7,
  337.2,
  336.6,
  336.4,
  336.3,
  335.9,
  335.1,
  335.1,
  333.6,
  328.9,
  326.1,
  324.4,
  324.9,
  326.2,
  327.9,
  328.9,
  329.3,
  329.5,
  328.9,
  328.7,
  329,
  329.2,
  329.5,
  329.8,
  330.4,
  328.8,
  327.6,
  333.1,
  334.6,
  335.4,
  336.5,
  335.8,
  335.9,
  336.7,
  336.7,
  338.4,
  338.4,
  339.5,
  347,
  340.5,
  338.2,
  337.9,
  337.9,
  337.4,
  337.8,
  338.2,
  338.5,
  338.5,
  338.7,
  338.8,
  338.7,
  338.2,
  337.8,
  337.1,
  336.5,
  335.5,
  335,
  334.5,
  333.8,
  333.1,
  330.6,
  327.9,
  326.6,
  325.4,
  324.7,
  323.5,
  322.7,
  321.9,
  322.1,
  322.1,
  322.4,
  322.9,
  323.1,
  323.5,
  324.7,
  326.6,
  328.7,
  331.4,
  332.2,
  340.7,
  345.2,
  347.7,
  347.6,
  344.1,
  341.8,
  338.8,
  354.8,
  338.2,
  330,
  331.2,
  331.1,
  323.5,
  325.9,
  324.5,
  324.9,
  322.8,
  317.8,
  302.3,
  277,
  247.3,
  265.8,
  292.4,
  311.8,
  282.7,
  254.8,
  264,
  298.8,
  311.6,
  316.6,
  316.8,
  322.1,
  323.9,
  319.8,
  318,
  318.3,
  311.9,
  307.2,
  301.6,
  264.1,
  298.7,
  306.8,
  299.1,
  261.6,
  282.9,
  309,
  316.7,
  318.1,
  318.6,
  319.7,
  320.9,
  320.8,
  320.6,
  319,
  320.5,
  329,
  322.5,
  320,
  308.5,
  252.6,
  241.5,
  263.9,
  279.9,
  300.3,
  285.2,
  284.2,
  280.8,
  279.9,
  279.6,
  280.3,
  281.8,
  283.4,
  287.2,
  289.5,
  291.7,
  293.6,
  293.6,
  292.8,
  298.6,
  302.5,
  288.7,
  296.7,
  315.3,
  301.4,
  271.1,
  292.8,
  287.8,
  305.9,
  294.1,
  274.3,
  277.9,
  304.2,
  290.9,
  279.9,
  302.5,
  333.9,
  322.5,
  321.8,
  316.8,
  315.8,
  315.2,
  340.7,
  308.4,
  330.5,
  292.2,
  282.9,
  284.5,
  283.1,
  302.8,
  345.1,
  345.5,
  345.6,
  315.2,
  340.5,
  322,
  288.5,
  296.9,
  338.9,
  307.5,
  322.1,
  295.6,
  272.9,
  282.8,
  337.9,
  311.3,
  286.4,
  271.8,
  265.6,
  273.3,
  321.4,
  280,
  273.7,
  314,
  329.9,
  329.5,
  318.2,
  291.5,
  331.5,
  321,
  333.4,
  343.1,
  339.9,
  336,
  274.3,
  329.6,
  343.2,
  339.3,
  341.6,
  329.4,
  281,
  265.5,
  286,
  274.3,
  269.6,
  274.3,
  281,
  282.9,
  281.4,
  280.3,
  285.9,
  293.2,
  294,
  303.5,
  308.8,
  314.9,
  320.7,
  324.9,
  325.8,
  330.7,
  336,
  341.1,
  339.2,
  336.2,
  339.5,
  341.2,
  337.7,
  337,
  337.2,
  338.2,
  338.7,
  339.5,
  337.1,
  336,
  335.4,
  335.6,
  335.4,
  334.5,
  328.2,
  329.7,
  339.2,
  347,
  347.2,
  354.3,
  358.9,
  360.7,
  362,
  366.9,
  367.8,
  352.5,
  375.1,
  284.4,
  259.2,
  283.7,
  306.7,
  301,
  306,
  291.9,
  283.6,
  285.5,
  287.1,
  295.1,
  297.1,
  297,
  297.6,
  299.8,
  299.2,
  297.5,
  301.2,
  301.9,
  305.6,
  301.8,
  301.5,
  302.6,
  301.5,
  306.4,
  304.8,
  305.4,
  304.1,
  300.2,
  301.1,
  304.1,
  305.6,
  308.3,
  310.5,
  309.6,
  303.6,
  288.5,
  269.5,
  258.2,
  261.5,
  258.7,
  281.1,
  294,
  269.7,
  269.7,
  265.4,
  266.2,
  326.9,
  282.1,
  249.1,
  254.5,
  286.9,
  289.5,
  276.5,
  294,
  298.3,
  284.7,
  306.4,
  311.2,
  312.1,
  313.4,
  314,
  314.2,
  313.4,
  314.2,
  316.2,
  317.2,
  317.4,
  316.9,
  318,
  317.5,
  317.2,
  317.5,
  317.9,
  318.4,
  319,
  318.9,
  318.5,
  320.5,
  319.9,
  319.2,
  317.4,
  317.5,
  317.6,
  317.3,
  317.5,
  317.6,
  317.2,
  317.1,
  317,
  317.4,
  316.3,
  315.7,
  314.7,
  313.1,
  320,
  314,
  289.4,
  232.5,
  237.8,
  237,
  235.3,
  233,
  240.9,
  247.2,
  251,
  255.1,
  256.3,
  257.7,
  258.9,
  261.5,
  262.7,
  263.8,
  265.5,
  267.1,
  268.3,
  282.3,
  295.1,
  296,
  283.9,
  274.2,
  280.2,
  271.7,
  265.9,
  266.6,
  266.4,
  266.9,
  267.5,
  265.6,
  265.5,
  264.8,
  274.4,
  276.1,
  276.9,
  271.1,
  277.2,
  262.2,
  251.4,
  281.2,
  284.6,
  293.9,
  295.8,
  294.9,
  285.4,
  259.8,
  230.4,
  231.9,
  251.7,
  259.3,
  236.1,
  235.7,
  237.6,
  238.8,
  242.7,
  245,
  266.5,
  290.1,
  307.7,
  312.1,
  310.6,
  310.8,
  310.5,
  309.9,
  310,
  309.3,
  310.8,
  312.2,
  313,
  314.2,
  314.6,
  316.4,
  316.1,
  317.8,
  318.9,
  320.1,
  320,
  321,
  321.1,
  322.2,
  324.5,
  326.8,
  329.6,
  332.8,
  333.8,
  335.2,
  335.6,
  336.2,
  335.7,
  334,
  333,
  332.9,
  346.5,
  340.1,
  326.8,
  328.5,
  329,
  329.9,
  331.9,
  332,
  329.8,
  330.6,
  331.4,
  331.8,
  331.6,
  332.2,
  331.8,
  331.1,
  330.2,
  329.6,
  329.5,
  329.2,
  329.1,
  329,
  329.1,
  329,
  329.2,
  329.3,
  329.5,
  329.2,
  328.8,
  328.9,
  328.5,
  327.9,
  326.8,
  325.8,
  326.2,
  327.3,
  328.8,
  330.4,
  332.2,
  332.8,
  333.9,
  334.9,
  332.7,
  330.3,
  329.1,
  328.7,
  328.4,
  328.2,
  348.7,
  336,
  327.9,
  327.6,
  327.5,
  327.3,
  325.7,
  325.1,
  324.7,
  324.5,
  326.1,
  326.6,
  327.3,
  326.6,
  326.7,
  326,
  325.4,
  324.1,
  321.1,
  321.8,
  319.2,
  316.2,
  319.7,
  319.7,
  319.8,
  320.3,
  321.6,
  324.3,
  324.9,
  325.2,
  325,
  324.8,
  324.4,
  323.1,
  326.8,
  327.7,
  327.5,
  327.4,
  328.8,
  329.3,
  329.6,
  329.2,
  327.8,
  326.1,
  325.1,
  323.1,
  321.8,
  321.7,
  332.9,
  326.3,
  322.6,
  321.9,
  322.1,
  322,
  322.1,
  321.7,
  321.4,
  321.7,
  321.7,
  321.7,
  321.7,
  321.3,
  321.7,
  321.4,
  321.3,
  321.9,
  321.3,
  317.3,
  315.7,
  317.9,
  316.6,
  312.8,
  277.8,
  248,
  247.3,
  246.8,
  247.7,
  273.9,
  257.8,
  272.3,
  313.2,
  321.1,
  326.1,
  326.6,
  327.8,
  329,
  330.3,
  332.2,
  333.9,
  336,
  340.1,
  342.5,
  342.2,
  342.6,
  341,
  341.5,
  340.2,
  345.4,
  336.6,
  332.6,
  331.3,
  330,
  328.7,
  327.9,
  327.6,
  325.3,
  317.1,
  316.1,
  315.2,
  316.1,
  316.5,
  316.9,
  316.2,
  315.8,
  315.5,
  316.1,
  314.6,
  314.5,
  316.4,
  314.4,
  314.3,
  314.4,
  314.2,
  315.5,
  315.7,
  314.5,
  314,
  313.4,
  313.3,
  311.8,
  311.1,
  309.6,
  308.5,
  308.6,
  308.1,
  308.5,
  308.6,
  309.4,
  308.4,
  304.7,
  285.4,
  281.1,
  290.9,
  293.8,
  303.8,
  319.1,
  308.1,
  301.7,
  295.1,
  301.2,
  301.3,
  295.3,
  294.4,
  277.4,
  232.9,
  231,
  229.1,
  229.4,
  230.4,
  231.3,
  231.3,
  232.3,
  241.6,
  234.9,
  230.4,
  232,
  231.2,
  228.5,
  228.8,
  234.1,
  237.8,
  233.9,
  235.2,
  253.6,
  283.7,
  243.7,
  237.2,
  236.2,
  238.9,
  240.4,
  238.1,
  251,
  261.5,
  257.8,
  254.5,
  238,
  251.7,
  276.3,
  301.2,
  263.7,
  301.3,
  309.6,
  311.9,
  317.9,
  313.5,
  314.2,
  314.3,
  314.9,
  315.5,
  315.7,
  316.5,
  317,
  317.5,
  317.8,
  318.5,
  319,
  319.7,
  319.9,
  319.9,
  320.4,
  320.5,
  320.9,
  321.1,
  321.3,
  321.4,
  321.6,
  321.6,
  321.7,
  322.3,
  322.8,
  321.9,
  321.5,
  320.4,
  320.3,
  319.8,
  320.1,
  320.7,
  321.7,
  323.4,
  325.4,
  327.3,
  329.2,
  328.4,
  328.1,
  328.2,
  326.6,
  323.7,
  322.7,
  322.2,
  321.9,
  321.8,
  338.7,
  325.8,
  322.7,
  321.8,
  320.1,
  319.8,
  318.9,
  318.2,
  317,
  317,
  316.1,
  317.2,
  318.3,
  319.4,
  316.7,
  307.2,
  311.3,
  311,
  313.6,
  313.8,
  308.5,
  304.2,
  306.6,
  313.1,
  315.2,
  317,
  316.6,
  317.3,
  309.7,
  308.5,
  302.5,
  302.3,
  313.2,
  321.5,
  324.6,
  326.5,
  327.6,
  328.7,
  329.4,
  330.2,
  330.6,
  331.7,
  333,
  334,
  335.2,
  337.1,
  338.3,
  338.8,
  343,
  341.3,
  341.2,
  342.2,
  342.5,
  342.9,
  343.6,
  343.6,
  344.5,
  344.8,
  345.3,
  345.8,
  345.1,
  344.9,
  345,
  344.4,
  344.2,
  344.3,
  336.3,
  329.2,
  329,
  330.3,
  331.5,
  330.8,
  329.5,
  326.4,
  328.4,
  330,
  329.8,
  328.8,
  326.7,
  326.7,
  326.8,
  324.4,
  320.9,
  325.2,
  334.5,
  339.1,
  312.9,
  282.9,
  266,
  280.7,
  293.9,
  296.3,
  313,
  312.5,
  316.3,
  318.7,
  334.3,
  301.9,
  253,
  266.8,
  269.4,
  252.8,
  284.7,
  293.6,
  296.9,
  243.4,
  249.2,
  266.4,
  279,
  287.7,
  291.2,
  297,
  297.6,
  299.6,
  305.1,
  309.1,
  308.5,
  318.7,
  323.6,
  326.1,
  326.9,
  326.8,
  326.7,
  326.6,
  325.7,
  325,
  324.5,
  324.4,
  324.3,
  324.4,
  325.3,
  327.1,
  327.7,
  329.3,
  328.4,
  311.5,
  305.9,
  310.1,
  303,
  310.1,
  310.8,
  313.8,
  329.4,
  326.3,
  356.2,
  312.3,
  332.9,
  322.1,
  309.8,
  306.9,
  302.3,
  270.3,
  263.7,
  266.3,
  276.7,
  299.1,
  306.4,
  315.3,
  325.6,
  330.1,
  330.4,
  330.8,
  331,
  329.8,
  330.3,
  330.5,
  331.6,
  332.1,
  331.6,
  333.5,
  333.4,
  335.3,
  337.5,
  338.7,
  341.8,
  338.3,
  337.4,
  335.6,
  326.1,
  322.3,
  339.5,
  329.2,
  315.7,
  279.2,
  301.5,
  321.2,
  346.7,
  349.1,
  347.8,
  346.7,
  346.7,
  349,
  361,
  355.8,
  352.4,
  351.3,
  350.9,
  351.2,
  349,
  347.1,
  347.2,
  345.8,
  345.1,
  344.9,
  344.6,
  343.5,
  341.3,
  338,
  335.7,
  332.3,
  330.3,
  328.4,
  326.2,
  323.9,
  320.6,
  318.1,
  316,
  315.2,
  315.3,
  315.6,
  314.2,
  316.7,
  312.9,
  310.8,
  309.3,
  310.4,
  312.4,
  311.4,
  318.7,
  319.3,
  324.2,
  336,
  334.5,
  342.6,
  348.8,
  345,
  283.8,
  264.8,
  270.8,
  266.5,
  313.7,
  293.7,
  264.9,
  255.5,
  265.2,
  285.1,
  301.2,
  307.1,
  308.7,
  306.7,
  318.8,
  331.7,
  334.3,
  337,
  339.1,
  339.3,
  340.8,
  341.7,
  343,
  343.9,
  344.3,
  343.7,
  343.2,
  342.5,
  341.1,
  333.4,
  326.4,
  334,
  322,
  301.9,
  276.9,
  258.1,
  262.6,
  260.7,
  257.4,
  279.4,
  315.8,
  341.9,
  351.7,
  349.7,
  342.6,
  331.2,
  314.5,
  325.1,
  341.1,
  345.9,
  350,
  351.8,
  364.3,
  355,
  350.9,
  349,
  348.2,
  346.3,
  334.4,
  327.6,
  330.7,
  334.2,
  311.2,
  315.6,
  339.6,
  322,
  337.5,
  324.9,
  316.6,
  306.9,
  312.6,
  319.9,
  314.9,
  331.8,
  308.4,
  295.8,
  300.5,
  287.3,
  290.4,
  314.6,
  272.5,
  277.8,
  289.6,
  326.9,
  335.5,
  338.2,
  328.7,
  339.2,
  336,
  338.1,
  339.9,
  338.5,
  343.6,
  345.9,
  346.5,
  345.7,
  347.8,
  348.6,
  350.7,
  351,
  358.2,
  355.5,
  354.7,
  356.7,
  357.6,
  354.7,
  338.2,
  272.2,
  260.6,
  256.2,
  254.5,
  249.9,
  246.4,
  243.9,
  243.1,
  244.6,
  245.6,
  245.8,
  245.8,
  244.4,
  243.3,
  242,
  240.6,
  239.6,
  238.4,
  238.6,
  240.4,
  242.8,
  242.4,
  242.4,
  246.9,
  250,
  243.2,
  245.6,
  249.5,
  260.4,
  277.9,
  299.8,
  283.7,
  316.7,
  337.2,
  335.2,
  327.2,
  336.6,
  332.5,
  325.7,
  324.6,
  313.7,
  344.3,
  327.8,
  308.3,
  308.7,
  297,
  297.2,
  310.1,
  317.3,
  323.5,
  321.3,
  329.1,
  328.2,
  334.4,
  338.4,
  339.9,
  340.4,
  340.8,
  340.9,
  342,
  343.1,
  345,
  348.1,
  351.3,
  355.2,
  359.5,
  361,
  361.6,
  360.9,
  361.4,
  359.9,
  359.5,
  359.2,
  358.5,
  358.1,
  359.2,
  358.4,
  359.7,
  359.7,
  359.5,
  361.4,
  361.8,
  362.4,
  363.3,
  363.6,
  362.6,
  362.8,
  364.4,
  364.8,
  373.6,
  365.4,
  361.7,
  361.7,
  362.2,
  363.5,
  361.7,
  361.3,
  360.7,
  359.3,
  359.5,
  359.6,
  359,
  359.9,
  361,
  359.8,
  359,
  358.9,
  359.5,
  358.5,
  359.1,
  357.6,
  353.5,
  348.1,
  337.3,
  331.3,
  324.7,
  335.3,
  295.4,
  319.1,
  330,
  341,
  342.5,
  336.6,
  335.7,
  326.8,
  320.5,
  314.9,
  320.8,
  329.7,
  325.5,
  328.1,
  332.4,
  332.7,
  331.9,
  333.1,
  332,
  334.9,
  343.8,
  336.7,
  333.6,
  332.3,
  331.7,
  331.8,
  331.7,
  330.7,
  329.5,
  327.4,
  326,
  325.4,
  325.2,
  324.1,
  321.9,
  320.7,
  317.1,
  303.2,
  290.9,
  249.1,
  245.7,
  260.2,
  270.9,
  254.6,
  244.4,
  240.6,
  239.2,
  239.1,
  239.3,
  238.2,
  237.2,
  236.3,
  234.1,
  236.2,
  237.9,
  239.4,
  240.7,
  241.8,
  242.8,
  245.6,
  269,
  266.2,
  303.1,
  295.7,
  290.7,
  269.2,
  249.9,
  271.9,
  315.5,
  267.7,
  243.6,
  245.7,
  248.2,
  251.1,
  252,
  249.1,
  245.6,
  250.5,
  248.6,
  248.2,
  245,
  245.6,
  311.2,
  305.7,
  314.5,
  311.1,
  307.4,
  303.3,
  270,
  275.3,
  312.8,
  311.6,
  310.3,
  281.7,
  262.9,
  271.3,
  278.1,
  276.6,
  274.2,
  281.4,
  305.1,
  301.6,
  255.6,
  242.5,
  244.3,
  248.5,
  265,
  263.3,
  289.3,
  274.8,
  304.9,
  313.7,
  303.4,
  301.9,
  279.7,
  275.6,
  338.6,
  282.1,
  251.2,
  265,
  274.2,
  284.4,
  275.1,
  286.9,
  317.9,
  296,
  279.7,
  298,
  313,
  315.3,
  308.8,
  303.2,
  272.7,
  275.6,
  272.1,
  252.9,
  263.5,
  278.6,
  312.3,
  313.8,
  314,
  308,
  303.9,
  314.6,
  318,
  312.2,
  306.7,
  284.8,
  276.6,
  271.9,
  260.6,
  279.5,
  301.1,
  292.5,
  300.5,
  304.2,
  285.3,
  285.9,
  284.9,
  282.2,
  279.9,
  284,
  285.3,
  285.4,
  282.9,
  299.7,
  285.3,
  277.7,
  280.9,
  275.2,
  252.6,
  246.2,
  251.5,
  247,
  263.7,
  262.7,
  254.4,
  271.8,
  302.8,
  299.6,
  312.5,
  324.7,
  329.5,
  323.7,
  321.8,
  323.4,
  324.3,
  324.8,
  328.3,
  328,
  330.2,
  331,
  332.1,
  332.7,
  332.1,
  332.4,
  333.7,
  334.3,
  334.9,
  336.1,
  337.2,
  338.3,
  340.5,
  341.7,
  342,
  335.1,
  339.7,
  338.7,
  308.7,
  315.4,
  322.5,
  298.6,
  326.7,
  346.1,
  329.9,
  322.8,
  312.3,
  305.6,
  307.8,
  318.8,
  329.1,
  329.3,
  330,
  339.7,
  328.3,
  332.7,
  342.7,
  351.1,
  352.7,
  349.9,
  349.5,
  349.2,
  348.6,
  350.7,
  352.1,
  352.3,
  352.8,
  353.5,
  353.3,
  353.9,
  354.7,
  354.8,
  354.1,
  355.2,
  356.9,
  358.9,
  358.2,
  332.9,
  315.9,
  329.5,
  327.6,
  348,
  330.6,
  323.1,
  320.3,
  320.1,
  318.3,
  316.5,
  322.9,
  333.9,
  284.6,
  331.2,
  263,
  255.1,
  250.7,
  272.8,
  276.4,
  316.3,
  306.4,
  317.7,
  326.1,
  285.5,
  272.7,
  250.4,
  245.6,
  246.2,
  245.5,
  274,
  314.3,
  321.4,
  321.2,
  320.2,
  310.8,
  305.8,
  315.9,
  304.7,
  244.6,
  241.3,
  241.4,
  237.9,
  235.9,
  235.1,
  246.4,
  239.8,
  263.8,
  243.5,
  243.2,
  262.4,
  286.2,
  301.2,
  307.3,
  312.8,
  322.2,
  326.5,
  323.6,
  320.7,
  326,
  316.3,
  323.5,
  336.8,
  331.1,
  326.6,
  328.8,
  332.5,
  335.1,
  336.3,
  335.1,
  337.5,
  340.3,
  342.2,
  343.1,
  345.7,
  348.4,
  348.7,
  331.5,
  339.3,
  292.5,
  329.4,
  312.2,
  293.7,
  251.6,
  247.9,
  247.7,
  247.5,
  249.6,
  251.7,
  252.3,
  265.1,
  248.4,
  246.4,
  245,
  245.3,
  249.1,
  253.2,
  257.6,
  263.1,
  286.9,
  292.8,
  296.2,
  304.8,
  308.5,
  311.1,
  319.6,
  316.8,
  322.7,
  323.6,
  324.8,
  355.4,
  346.8,
  340,
  346.5,
  346.1,
  336.8,
  330.2,
  341.5,
  331.3,
  335.2,
  330.4,
  340.4,
  345.5,
  346.2,
  345.4,
  346.7,
  345.5,
  344.7,
  344.9,
  340.7,
  345.9,
  348.4,
  348.8,
  348,
  346,
  348.5,
  349.2,
  350.3,
  350,
  351.2,
  351,
  351.1,
  351.9,
  353,
  353.5,
  354.7,
  355.4,
  357.8,
  356.7,
  356.5,
  357,
  357.2,
  357.9,
  357,
  354.2,
  352.9,
  349.4,
  354.2,
  358.1,
  323.9,
  282.7,
  312.5,
  336.2,
  335,
  339.3,
  337.3,
  326.8,
  322.6,
  322.4,
  333.3,
  344.4,
  331.6,
  336.4,
  322.3,
  315,
  281.4,
  310.3,
  310.3,
  312.4,
  327.1,
  339.6,
  342,
  337.4,
  345.6,
  343.2,
  334.2,
  345.3,
  346.9,
  348.3,
  349.4,
  350.2,
  351.6,
  353.4,
  355.3,
  356.6,
  357.7,
  358.9,
  359.6,
  359.5,
  359,
  353.5,
  353.2,
  351.4,
  352.3,
  353,
  353.9,
  362.5,
  353,
  349.7,
  352.2,
  351.8,
  354.1,
  352,
  348.3,
  324.2,
  344.5,
  352.2,
  350.8,
  350.9,
  350.9,
  351,
  350.3,
  340.6,
  337.2,
  333.9,
  295.5,
  290.5,
  288.2,
  321.5,
  305.1,
  288.7,
  290,
  292.1,
  308.8,
  312.8,
  334.4,
  333.6,
  336.2,
  337.9,
  331.3,
  326.6,
  309.8,
  290,
  292.6,
  310.8,
  306.6,
  313.2,
  324.2,
  330.9,
  346.7,
  346.5,
  340.4,
  348.4,
  353.6,
  362.8,
  357.1,
  352.4,
  352.6,
  350.3,
  351.1,
  349,
  347.1,
  345.1,
  345.3,
  341.2,
  340.8,
  338.9,
  341.9,
  331.5,
  316.3,
  309.8,
  307.3,
  317.2,
  330.7,
  330.7,
  288.6,
  315.6,
  334.3,
  351.2,
  350.5,
  359.6,
  357.3,
  356.3,
  354.6,
  358.3,
  359.6,
  348.9,
  343.4,
  346.1,
  350.9,
  348.6,
  352.1,
  343.7,
  340.5,
  341.1,
  343.2,
  335.4,
  345.1,
  344.1,
  341.9,
  273.7,
  330.8,
  346.2,
  289.8,
  281,
  293.2,
  311.1,
  321,
  334.1,
  346.5,
  349.3,
  351.3,
  353.4,
  355.3,
  360.7,
  362.9,
  364,
  364.1,
  365.3,
  366.6,
  364.3,
  344.4,
  348.8,
  326.8,
  330,
  349.3,
  346,
  322.5,
  338.3,
  344.4,
  346.6,
  318.8,
  327.8,
  339,
  340,
  346.3,
  332.4,
  326.1,
  328.3,
  303.2,
  332.4,
  301.8,
  316.7,
  342.5,
  326.3,
  322.1,
  326,
  329.5,
  331.5,
  337,
  353.1,
  306.8,
  287.8,
  284.8,
  289,
  294,
  339,
  350.7,
  351.6,
  351.5,
  359,
  352.2,
  342.9,
  347.8,
  337.6,
  349.3,
  348.7,
  352.4,
  345.9,
  326.6,
  344.1,
  341.3,
  336.2,
  331.4,
  313,
  306.7,
  315.7,
  267.7,
  271.5,
  279.1,
  288.6,
  300.3,
  326,
  328.1,
  336.8,
  335.1,
  342.1,
  339.6,
  338.7,
  337.7,
  343.4,
  341.5,
  338.8,
  339.5,
  336.6,
  338.5,
  325.2,
  330.6,
  345.3,
  342.1,
  335.9,
  334.6,
  319.4,
  334.8,
  338.9,
  338.6,
  329.7,
  337,
  339,
  340.8,
  341.2,
  338.4,
  336.9,
  336.1,
  336.6,
  332.9,
  332.5,
  330.9,
  323.4,
  286.1,
  247.7,
  293.1,
  298.5,
  246.9,
  252.9,
  269.4,
  279.9,
  284.6,
  283.3,
  272.3,
  249.3,
  307.2,
  329.2,
  341.9,
  341.7,
  322.8,
  325.6,
  326.4,
  330,
  322,
  324.8,
  324.9,
  328,
  316.5,
  305.2,
  301.1,
  354,
  314.6,
  303.3,
  318.3,
  326.9,
  324.9,
  325.3,
  323.4,
  307.9,
  320,
  314,
  301.4,
  285,
  293.1,
  291.3,
  281.8,
  278.8,
  275,
  267.8,
  269,
  268.9,
  264.4,
  266.7,
  269.4,
  267.8,
  266.1,
  265.2,
  270,
  270.5,
  274.6,
  271.1,
  265.5,
  268.4,
  272.8,
  283.3,
  292.8,
  295.1,
  291.4,
  291.6,
  285.4,
  293.7,
  307.4,
  310.6,
  319.2,
  317,
  315.6,
  314.6,
  316,
  359.2,
  328.6,
  312.7,
  304.7,
  297.1,
  306.1,
  293,
  334.5,
  340.8,
  349.8,
  352.6,
  357.9,
  355.3,
  356.8,
  358.6,
  359.5,
  359.3,
  358.9,
  357.4,
  350.2,
  327.6,
  307.7,
  281.7,
  279.2,
  287.7,
  297.4,
  305,
  309.3,
  312.1,
  308.9,
  305.3,
  315.5,
  290.3,
  248.6,
  255.2,
  259.6,
  265,
  270.1,
  273,
  279.5,
  288.1,
  294.6,
  302.9,
  301,
  281.8,
  278.7,
  281.5,
  282,
  347,
  347.6,
  352.2,
  334.9,
  303.7,
  317.6,
  342.2,
  353,
  350.9,
  358.3,
  361.4,
  359.1,
  357.3,
  334.1,
  338,
  347.2,
  346.5,
  360.1,
  360.3,
  360.6,
  361.3,
  361.9,
  361.1,
  361.3,
  361.1,
  360.5,
  360.6,
  359.7,
  359.7,
  360.2,
  360,
  360.5,
  360.3,
  361.2,
  361.5,
  360.8,
  347.8,
  339.6,
  364.4,
  364.5,
  364.6,
  363.6,
  363.7,
  365.5,
  369.1,
  353.7,
  347.2,
  345.8,
  363.1,
  350.9,
  308.5,
  270.7,
  272.3,
  282.9,
  278.7,
  269.7,
  268.3,
  279.3,
  301.7,
  292.4,
  286.3,
  289.5,
  295.3,
  301.3,
  303.3,
  298.6,
  294,
  300.9,
  288.2,
  284.9,
  273.8,
  266.8,
  265.5,
  264.3,
  262.4,
  291.8,
  290.4,
  262,
  257.4,
  263.6,
  281.4,
  255.1,
  252.3,
  250.5,
  253,
  256.3,
  259.3,
  260.7,
  273.8,
  270.2,
  268.6,
  274.3,
  292.6,
  300.3,
  299.5,
  307.7,
  351,
  328.1,
  316.2,
  321.7,
  324.3,
  322,
  324.5,
  323.7,
  323.1,
  315.5,
  321.4,
  324.1,
  317.4,
  314.5,
  307.2,
  304.1,
  296.9,
  279.1,
  318.1,
  276.7,
  269,
  273.6,
  274.6,
  274.1,
  273.9,
  270.7,
  265.6,
  262.3,
  260.8,
  254.9,
  250.5,
  251.9,
  256.7,
  261.3,
  266.3,
  272.7,
  306.1,
  327.1,
  334.6,
  339.5,
  339.4,
  339.5,
  337.3,
  318.7,
  311.7,
  325.2,
  311.7,
  315.3,
  327.9,
  334.9,
  312.6,
  304.9,
  302.4,
  321.9,
  327.5,
  322,
  307.9,
  307.6,
  318.7,
  304.9,
  301,
  300.2,
  313.5,
  314.1,
  298.3,
  294.6,
  293.5,
  293.6,
  292.8,
  290.1,
  289.5,
  288.8,
  289.1,
  291.2,
  295.3,
  297.5,
  321.1,
  355.6,
  358.6,
  357.5,
  357.1,
  354.4,
  342.4,
  345,
  355.5,
  356.4,
  314,
  349.5,
  348.5,
  341.7,
  299.3,
  283.4,
  283.9,
  285.8,
  279.5,
  277.6,
  277.5,
  311.5,
  282.1,
  295.1,
  340.7,
  342.9,
  326.8,
  329,
  343.9,
  337.9,
  307.5,
  263.5,
  262.8,
  261.8,
  265.8,
  307.8,
  329.9,
  339.7,
  344.3,
  344.7,
  344.7,
  345,
  347.2,
  347.8,
  348,
  348.3,
  348.6,
  349,
  349.3,
  350.5,
  351.1,
  350.8,
  350.9,
  353.2,
  360,
  317.9,
  272.8,
  295.2,
  310.5,
  312.2,
  303.6,
  286.3,
  280.6,
  306.8,
  296.4,
  298.7,
  322.7,
  284.3,
  276.9,
  314.1,
  275.6,
  267.1,
  264,
  263,
  262.3,
  259.8,
  269.7,
  276.2,
  258.5,
  259,
  258.7,
  263.2,
  269,
  263.2,
  260.5,
  257.5,
  257.3,
  285.9,
  260.4,
  264.1,
  330.7,
  338,
  338.2,
  338,
  338.6,
  340.3,
  339.4,
  337.3,
  334.7,
  319.6,
  279.9,
  291.4,
  306.3,
  301.5,
  308.1,
  301.8,
  298.5,
  302.8,
  306.3,
  310.3,
  330.6,
  355.7,
  348.6,
  336.5,
  328.6,
  336,
  341.6,
  358.1,
  339.3,
  334.6,
  324.4,
  316.3,
  315.9,
  305.1,
  306.4,
  308.9,
  303.6,
  320.3,
  324.2,
  308.5,
  310.3,
  318.8,
  320.5,
  301.9,
  323.6,
  327.3,
  325,
  325.2,
  296.5,
  297.7,
  303.1,
  290.8,
  318.8,
  336.6,
  327.6,
  340.1,
  310.3,
  282.5,
  318,
  344.8,
  349.3,
  351.3,
  353.3,
  354.3,
  356.8,
  359,
  349.4,
  350.3,
  362.6,
  355.4,
  348.9,
  352.7,
  337.8,
  321.3,
  292.8,
  328.3,
  297.8,
  290.3,
  289.2,
  287,
  285.5,
  285,
  284.1,
  282.4,
  282.8,
  285.3,
  285.5,
  281.6,
  280.1,
  280.4,
  293.6,
  315.8,
  332.2,
  342.2,
  347.7,
  349.1,
  348.7,
  346.7,
  345.8,
  345.2,
  345.1,
  343.4,
  342.4,
  340.5,
  336.7,
  331.2,
  324,
  315.4,
  328.3,
  324.3,
  313,
  282.2,
  270.3,
  268.6,
  276.4,
  279.4,
  281.7,
  282.2,
  282.2,
  282.5,
  284.5,
  284.7,
  282.9,
  329.7,
  292.9,
  281.8,
  281.6,
  280.4,
  277.6,
  276.1,
  274.5,
  273.4,
  270.8,
  270.2,
  269.5,
  268.4,
  268.2,
  267,
  268.5,
  268.6,
  268.7,
  268.3,
  267.2,
  267.1,
  264.4,
  262.9,
  261.5,
  263.3,
  263.2,
  264.1,
  261.9,
  255.7,
  254.1,
  258.9,
  259.8,
  265,
  271,
  276,
  279,
  282.3,
  282.8,
  276.6,
  286.2,
  289.2,
  289.4,
  288.8,
  288.4,
  289.2,
  286.6,
  288.5,
  290,
  345.3,
  307,
  293.1,
  287,
  282.9,
  282.2,
  282.4,
  280,
  272.5,
  313.1,
  338.6,
  338.1,
  337,
  336.9,
  334.6,
  334.6,
  334.3,
  333.4,
  333.6,
  333.2,
  333.2,
  332.9,
  333.6,
  334,
  334.3,
  332.9,
  331.6,
  332,
  332.4,
  332.6,
  332.2,
  331.9,
  333.5,
  334.8,
  336.3,
  336.4,
  337.7,
  338.7,
  335.9,
  300,
  277.4,
  278.1,
  278.6,
  279.1,
  275.4,
  271.5,
  269.5,
  268.6,
  316.4,
  281.5,
  271.3,
  272.7,
  273,
  273.5,
  271.1,
  268.4,
  267.2,
  267,
  298.1,
  317.7,
  315.9,
  312.9,
  320.3,
  320.8,
  324.8,
  318.9,
  327.4,
  329.7,
  327.5,
  327.9,
  325.4,
  321.5,
  316.9,
  323.1,
  325.3,
  324.4,
  326.4,
  326.1,
  323.4,
  323.9,
  324.6,
  326.3,
  301.6,
  265.5,
  264.7,
  269,
  266.1,
  274.3,
  275.7,
  278,
  280.3,
  280.2,
  286.2,
  292,
  283,
  283.8,
  331.8,
  298.6,
  287.9,
  287,
  290.5,
  289.9,
  286.4,
  284.3,
  280.2,
  277.9,
  280.1,
  285.9,
  292.6,
  338.9,
  295.5,
  277.3,
  277.3,
  285.1,
  338.5,
  345.3,
  345.1,
  344.7,
  347.5,
  345.8,
  342,
  298.3,
  279.5,
  274.1,
  271.1,
  268.7,
  267.5,
  269.4,
  271.8,
  276.3,
  280.7,
  283.7,
  286,
  288.3,
  291.2,
  317.3,
  331.7,
  337.2,
  326.9,
  323,
  332.3,
  320.3,
  332.9,
  325.4,
  359.1,
  340.1,
  315.7,
  342.4,
  350.6,
  348.7,
  345.6,
  345.1,
  344.7,
  344.9,
  345.1,
  345.5,
  346.6,
  346.2,
  345.8,
  344,
  338.7,
  342.3,
  341.8,
  335.2,
  336.4,
  335.7,
  336.9,
  335.9,
  338.5,
  342.3,
  343.9,
  340.4,
  345.1,
  347.2,
  348.4,
  349.6,
  350.8,
  351.8,
  352.2,
  355.6,
  357.7,
  358.7,
  360.3,
  361.7,
  362.4,
  363,
  363.2,
  364.1,
  362.9,
  361.7,
  361.4,
  362.1,
  388.9,
  368.4,
  359.7,
  356.2,
  353.6,
  344.7,
  307.1,
  342.7,
  324.7,
  339.7,
  344,
  348.3,
  342.7,
  334.1,
  338,
  338.3,
  315,
  342.8,
  343.2,
  341.5,
  342.7,
  340.5,
  342.6,
  343.8,
  342.6,
  343.3,
  343,
  344.8,
  346.2,
  332.8,
  319.8,
  332.1,
  351.2,
  351.8,
  351.5,
  354.3,
  356,
  359.6,
  359.4,
  359.9,
  361.2,
  362.7,
  363.3,
  364,
  363.6,
  363.5,
  364.8,
  364.7,
  367,
  364.6,
  362.9,
  362.7,
  363.1,
  362.8,
  362.9,
  362.3,
  361.3,
  359.6,
  360.5,
  360.1,
  357.7,
  356.9,
  355.9,
  355.7,
  355.6,
  354.1,
  352.9,
  352.5,
  352.6,
  352.4,
  352.3,
  353,
  353.1,
  353.4,
  354.1,
  354.9,
  356.1,
  356.9,
  357.9,
  359.1,
  360.5,
  363.6,
  365.6,
  365.9,
  365.3,
  364.9,
  364.7,
  364.6,
  365.2,
  365.2,
  365,
  365.7,
  364.6,
  364.2,
  363.1,
  355.4,
  366.2,
  356.3,
  350.4,
  352.5,
  352.9,
  353.9,
  354.4,
  355.3,
  353.6,
  353.2,
  355.5,
  355.4,
  355.6,
  356.8,
  357.9,
  358.1,
  359.5,
  358.7,
  357.9,
  356.8,
  355.8,
  354.7,
  353.2,
  346.5,
  348.3,
  344.1,
  340.1,
  347.4,
  342,
  293,
  311.6,
  334.7,
  343.1,
  342.9,
  346,
  346.3,
  342.1,
  346.4,
  322.7,
  340.9,
  341.3,
  339.1,
  337.6,
  339.2,
  349,
  344.3,
  340.9,
  336.2,
  369.2,
  340.4,
  329.9,
  335.7,
  333.1,
  332.5,
  321.5,
  321.1,
  290,
  276.3,
  275.1,
  265.8,
  261.8,
  261.9,
  259.6,
  261.9,
  262.5,
  314.6,
  328.5,
  308.4,
  299.7,
  331.1,
  336.1,
  338,
  339.7,
  339.4,
  337.4,
  337.9,
  334.6,
  332,
  346.8,
  348.8,
  349.3,
  351.5,
  354.5,
  354.8,
  356.5,
  357.1,
  358.7,
  354.7,
  353.3,
  352.8,
  348.7,
  345.3,
  346.1,
  346.4,
  349.5,
  350.8,
  355.2,
  354.2,
  349.7,
  338.8,
  340.2,
  336.8,
  334.5,
  301.7,
  302.5,
  296.1,
  317.5,
  341.3,
  333,
  326.9,
  326.9,
  330.4,
  337.9,
  339.3,
  337.6,
  337.5,
  339.7,
  344,
  343.5,
  344.3,
  345.2,
  344.9,
  345.2,
  344.3,
  345.1,
  345.3,
  334.5,
  342.4,
  344.3,
  343,
  343.7,
  340.3,
  339.1,
  352.9,
  359.4,
  355.7,
  332.5,
  332.5,
  331.7,
  335.8,
  335,
  332.2,
  332.1,
  326.8,
  332.9,
  325.6,
  321.8,
  321,
  319.3,
  317,
  316.6,
  315.5,
  316.2,
  316.4,
  316.9,
  315.9,
  313.7,
  312.7,
  310.7,
  311.1,
  310.1,
  309.7,
  308.5,
  308.5,
  308.2,
  307.3,
  306.9,
  307,
  305.1,
  304.5,
  307,
  270.5,
  237.6,
  249.4,
  301.3,
  309.2,
  309.4,
  305.9,
  305.6,
  314,
  312.3,
  317.2,
  322.4,
  324.1,
  326.1,
  325.1,
  328.3,
  329.9,
  327.2,
  332.4,
  337.6,
  339.4,
  355.5,
  367.4,
  343.7,
  341.2,
  341.2,
  340.7,
  340.8,
  341,
  340.9,
  341,
  341.3,
  339.7,
  338.7,
  337.9,
  337.4,
  336.9,
  336.8,
  337.2,
  337.1,
  331,
  267.3,
  294.5,
  298.5,
  309.7,
  329.4,
  329.6,
  317.5,
  323.6,
  316.8,
  329.7,
  325.3,
  322.8,
  309.3,
  324.7,
  320.6,
  315.9,
  311.5,
  331.5,
  318.5,
  323.4,
  331.8,
  318.5,
  299,
  298.9,
  311.6,
  280.3,
  266.6,
  316.2,
  290.9,
  316.7,
  319.7,
  290,
  261.1,
  290.1,
  265.1,
  234.9,
  236.6,
  239.5,
  242.3,
  242.9,
  242.4,
  242.5,
  243.1,
  240.8,
  242.4,
  244.3,
  244.1,
  244.4,
  244.4,
  250,
  252.7,
  245.2,
  250.9,
  248.9,
  240.6,
  240.9,
  233.9,
  249.4,
  279.4,
  262.4,
  305.8,
  309.4,
  312.9,
  318,
  312.4,
  304.9,
  265.9,
  265.5,
  268.9,
  268.9,
  276.7,
  265.3,
  260.6,
  258,
  263.8,
  267.3,
  281.8,
  306.7,
  298.2,
  310.5,
  326,
  317.7,
  322.4,
  321,
  318.2,
  314.9,
  296.9,
  318.5,
  325.4,
  322.8,
  324.1,
  327.9,
  325.5,
  322,
  319.7,
  318.2,
  306.4,
  304.1,
  310.1,
  320.9,
  320.7,
  318.5,
  320,
  332.7,
  335,
  335.4,
  335.6,
  335.3,
  331.6,
  336.2,
  337.3,
  338.8,
  339.2,
  340.4,
  342,
  342,
  339.9,
  336.6,
  337.1,
  337.5,
  339.8,
  344.9,
  344.6,
  345.1,
  345.3,
  350.8,
  348.5,
  345.4,
  344.7,
  344.3,
  345.2,
  345.1,
  345.5,
  345,
  343.2,
  343.2,
  343,
  343.5,
  343.2,
  341.7,
  341,
  340.8,
  341.1,
  341.1,
  341.1,
  340.6,
  340,
  339.7,
  338.3,
  337.5,
  337.7,
  338.9,
  340.6,
  342.9,
  344.2,
  344.6,
  346.6,
  350.6,
  353.1,
  357.3,
  357.9,
  346.2,
  340.3,
  341.8,
  341.1,
  337.1,
  336.7,
  335,
  333.2,
  332.1,
  329.4,
  330.9,
  334.2,
  344.5,
  346.4,
  346.4,
  346.5,
  345.4,
  346,
  344.7,
  345.1,
  346.3,
  346.8,
  346.2,
  346,
  346.3,
  346.6,
  346.6,
  346.6,
  346.3,
  346.3,
  345.1,
  344.5,
  344.2,
  344.3,
  344.1,
  343.4,
  343.5,
  343.2,
  343.5,
  344.3,
  344.9,
  347.2,
  353.2,
  361,
  369.1,
  364.6,
  367.8,
  372.1,
  376.7,
  359.2,
  339.2,
  341.6,
  341.5,
  343.1,
  339.6,
  341.7,
  342.9,
  340.4,
  338.4,
  338,
  356.4,
  338.4,
  299,
  285.6,
  296.1,
  313.1,
  322.7,
  296.7,
  293.9,
  285,
  284.7,
  285.7,
  291.3,
  284.8,
  282.4,
  290.9,
  282,
  309.7,
  325,
  325.9,
  329.2,
  332.6,
  331.2,
  328.8,
  329,
  329.6,
  329.2,
  323,
  319.8,
  324.9,
  334.1,
  335.8,
  335.3,
  329.2,
  343.2,
  353.9,
  354.7,
  353.2,
  351.3,
  350.5,
  356.7,
  356.2,
  352.9,
  352.1,
  359.7,
  359.9,
  360.5,
  361.6,
  375.6,
  365.7,
  362,
  364,
  362,
  363,
  363.4,
  364.2,
  364.6,
  365,
  365.2,
  365.8,
  366.4,
  365.3,
  355.9,
  352.8,
  330.1,
  319.9,
  305.1,
  327.3,
  299.2,
  289,
  281.9,
  274,
  272.9,
  276.2,
  273.9,
  269.3,
  267.1,
  267,
  268.1,
  282.4,
  295.6,
  293.8,
  334.4,
  337,
  339.2,
  334.1,
  336.5,
  335.2,
  308.6,
  329,
  293.3,
  334.7,
  319.3,
  295.8,
  326.1,
  343,
  366.4,
  356.8,
  352.1,
  345.1,
  347.2,
  357.3,
  359.7,
  361.2,
  361.1,
  361.8,
  363.4,
  361.5,
  360.7,
  360.4,
  360.7,
  360.5,
  348.3,
  338.6,
  337.2,
  333.5,
  319,
  327.8,
  329.3,
  329,
  330.6,
  329.7,
  331.9,
  330.6,
  329.5,
  327.6,
  320,
  320.2,
  314.4,
  318.8,
  317,
  310.6,
  311,
  322.2,
  326,
  331.9,
  329.1,
  326.5,
  324.5,
  322.5,
  320,
  320,
  291.2,
  317.5,
  343.4,
  329.1,
  327.4,
  329,
  326.6,
  325,
  318.1,
  285.5,
  257.2,
  298.3,
  279.8,
  287.1,
  265.9,
  251.9,
  263.2,
  256.2,
  249.1,
  248,
  250.5,
  254,
  254.4,
  261.2,
  291.2,
  317.2,
  320.2,
  287.7,
  276.8,
  314,
  317.4,
  323.4,
  307.5,
  294.8,
  299.6,
  301,
  318.3,
  329.2,
  308.1,
  330.3,
  328.7,
  322.3,
  335.4,
  335.3,
  326.8,
  326,
  335.9,
  331.5,
  315.2,
  333.6,
  358.6,
  335.2,
  306.7,
  310.7,
  328.7,
  336.1,
  336,
  336.6,
  336.1,
  336.4,
  317,
  300.6,
  334.9,
  333.9,
  306.3,
  269.6,
  263.7,
  282.7,
  305.7,
  300.9,
  290,
  268.5,
  301.2,
  323.9,
  285.8,
  302.9,
  311.8,
  265.3,
  258.5,
  262.5,
  275.5,
  277.2,
  319,
  319.9,
  293,
  285,
  290.4,
  295.5,
  339,
  346,
  342.1,
  333.1,
  332.7,
  334.9,
  291.4,
  282.9,
  280.3,
  279.4,
  356.3,
  296.8,
  271.8,
  271.8,
  269.2,
  270,
  269.4,
  270.4,
  269.5,
  268,
  267.7,
  266.9,
  268.5,
  268.2,
  270.1,
  275,
  269.9,
  275.5,
  268.3,
  266.8,
  267.2,
  272.6,
  277.5,
  279.2,
  277.7,
  283.1,
  266.7,
  254.7,
  237.6,
  248.4,
  266.6,
  271.7,
  275.2,
  278.8,
  282,
  283.9,
  283.3,
  279.3,
  287.9,
  289.4,
  292.9,
  290.6,
  286.8,
  285.7,
  283.8,
  281.9,
  279.5,
  277.9,
  351.4,
  302.3,
  277.2,
  277.4,
  276.8,
  281.7,
  286.5,
  286.4,
  284.9,
  285.1,
  286.2,
  283.5,
  278.7,
  279.4,
  275.6,
  273.4,
  273.4,
  273.8,
  273,
  276.6,
  273.4,
  271.7,
  274.4,
  275.2,
  276.3,
  273.8,
  265.7,
  259.6,
  261.7,
  266,
  270.8,
  275.6,
  278.6,
  282.1,
  285,
  287,
  286.6,
  281.9,
  291.4,
  293.4,
  294.6,
  294,
  293.6,
  293.2,
  290.9,
  289.4,
  285.4,
  282.7,
  360.2,
  307.1,
  277.3,
  277.9,
  276.3,
  272.9,
  271.7,
  270.5,
  267.7,
  273.5,
  276.3,
  274.8,
  274.8,
  276.8,
  279.5,
  282.2,
  279,
  279.6,
  278.8,
  278.7,
  280.1,
  277.5,
  275.8,
  310.6,
  331.1,
  330.3,
  327.8,
  328.5,
  331,
  334.7,
  337.1,
  340.1,
  344.2,
  345.5,
  347.9,
  347.3,
  348.9,
  348.4,
  347.9,
  342.5,
  347.5,
  351.7,
  351.1,
  349.4,
  335.8,
  328.2,
  336.2,
  305.5,
  325.2,
  351.9,
  342.1,
  312.8,
  304.2,
  309.7,
  289.5,
  292.2,
  325.2,
  343.9,
  338.7,
  336.1,
  337.4,
  338,
  340.7,
  339.7,
  341.3,
  344,
  345,
  344.8,
  338,
  338.7,
  339.5,
  333.8,
  312.9,
  329.6,
  339,
  340.2,
  334.6,
  288.5,
  311.5,
  344.3,
  344.1,
  344.5,
  334.7,
  335.2,
  346.3,
  344.9,
  346.8,
  345.3,
  339.3,
  338.3,
  317.7,
  299.6,
  292.8,
  271,
  270.5,
  274.8,
  337,
  313.2,
  328.5,
  273.5,
  250.4,
  250.3,
  251.7,
  252.9,
  251.7,
  253.4,
  253.4,
  252.3,
  251.8,
  264.7,
  273.6,
  283.2,
  275,
  251.3,
  277,
  249.2,
  243.6,
  238,
  242.7,
  280.1,
  263.4,
  304,
  304,
  310.6,
  270.1,
  316.7,
  280.5,
  332.3,
  332.2,
  301.3,
  305.7,
  289.5,
  321.9,
  302,
  297,
  296.3,
  309,
  310.5,
  303.9,
  296.9,
  278.3,
  268.7,
  307.7,
  281.2,
  342.6,
  314.3,
  273.9,
  276.9,
  310.1,
  291.8,
  291.8,
  293.4,
  295.9,
  305.7,
  312.8,
  314.7,
  317.5,
  319.8,
  321.6,
  325.9,
  327.8,
  329.1,
  332.2,
  334.9,
  337,
  338.8,
  342.4,
  346.6,
  350.3,
  353.3,
  354.9,
  355.1,
  354.5,
  355,
  355.4,
  356.5,
  356,
  356.6,
  356.6,
  356.4,
  356.2,
  357.9,
  359.2,
  357.9,
  359.5,
  360.2,
  360.2,
  359.9,
  359.9,
  358.6,
  358.5,
  360.5,
  370.7,
  366.6,
  361.5,
  361,
  361.6,
  362.2,
  354,
  290.3,
  338.1,
  330.9,
  334.8,
  336.2,
  330.4,
  325.1,
  323.4,
  321.2,
  319.1,
  317.1,
  313.4,
  301,
  252.6,
  251.4,
  262.7,
  290.7,
  248.7,
  244.1,
  239.7,
  234.7,
  238.7,
  250.4,
  264.2,
  264.3,
  261.8,
  285.3,
  274.6,
  282.8,
  282.1,
  281.6,
  306.4,
  294.3,
  313.5,
  294.8,
  289.6,
  287.7,
  272.1,
  262.4,
  274.1,
  309.8,
  292.1,
  287.6,
  257.6,
  244,
  246.2,
  241.3,
  238.2,
  237.9,
  239.8,
  239.4,
  236.1,
  236.6,
  235.6,
  237.3,
  236.5,
  237.3,
  239.1,
  239.4,
  238,
  239.4,
  243.3,
  238.8,
  238.2,
  240.9,
  241.5,
  238.1,
  232.9,
  231.8,
  234.6,
  237.2,
  239.7,
  243.8,
  248.3,
  249.7,
  254.2,
  253.2,
  270.8,
  262.1,
  287.3,
  290.1,
  259.1,
  259.6,
  259.7,
  258.7,
  257.7,
  256.4,
  255.2,
  254.5,
  365.5,
  301.4,
  265.6,
  263.7,
  263.5,
  261.4,
  261.5,
  259.6,
  257.6,
  258.1,
  259.1,
  260.8,
  257.9,
  256.3,
  257.3,
  255.8,
  253.1,
  252.7,
  251.6,
  250.1,
  252.1,
  252.6,
  251.3,
  252.2,
  245,
  239.9,
  242,
  244.8,
  248.9,
  256.6,
  262.6,
  263.3,
  266.1,
  268.8,
  272.5,
  275.7,
  276.1,
  272.5,
  274.6,
  277.9,
  279.2,
  279.9,
  280.1,
  280.1,
  278.1,
  275.9,
  274.9,
  275.6,
  276.2,
  305.9,
  286.3,
  285.6,
  282.8,
  282.5,
  279.1,
  275.6,
  274,
  281.6,
  292.3,
  302.3,
  299.2,
  290.2,
  294.6,
  288.3,
  280.1,
  294.4,
  294.7,
  296.6,
  291.9,
  292.7,
  289.8,
  287.5,
  295.6,
  305.7,
  292.1,
  296.1,
  303.6,
  311.3,
  309.9,
  303.8,
  301.3,
  307.6,
  315.9,
  321.7,
  320.4,
  322,
  320.9,
  317,
  307,
  310.9,
  310.1,
  307.4,
  301.1,
  293.7,
  291.3,
  287.4,
  286.8,
  328.5,
  292.3,
  283.1,
  282.1,
  284.3,
  278.1,
  280.8,
  281.2,
  278.4,
  277.8,
  274.9,
  272.2,
  270.7,
  270.4,
  272.9,
  276.1,
  277.7,
  279,
  290.1,
  289,
  284.2,
  282.7,
  289.8,
  280.1,
  291.5,
  317.3,
  308.3,
  326.6,
  309.1,
  266.6,
  274.9,
  281.1,
  288.3,
  292,
  295.8,
  295,
  293.1,
  300.5,
  302.5,
  304,
  305.6,
  310.5,
  311.5,
  303.6,
  300.7,
  299.6,
  299.6,
  298.2,
  344.2,
  302.6,
  289.3,
  287.6,
  285.1,
  286.3,
  284.9,
  281.1,
  282.2,
  278.3,
  277.7,
  278.3,
  274.9,
  277.3,
  276.5,
  277,
  276.7,
  276.7,
  303.8,
  338.6,
  343.2,
  343.2,
  342.3,
  345.9,
  344.4,
  337.5,
  344.6,
  344.8,
  315.3,
  342,
  347.5,
  346.1,
  341.6,
  346.6,
  339.1,
  334.4,
  322,
  318.5,
  322,
  297.7,
  311.7,
  303.5,
  295.2,
  301.5,
  316.5,
  304.1,
  292,
  300.2,
  336.2,
  324.5,
  300,
  298.6,
  298.8,
  311.6,
  301,
  268,
  250.9,
  263.2,
  298,
  286.1,
  260.6,
  262.3,
  313.9,
  306.3,
  302.9,
  288.6,
  331.6,
  318.5,
  308.3,
  302.2,
  324.8,
  312.4,
  273.2,
  295.6,
  281.8,
  309.3,
  318.3,
  313.7,
  306.7,
  314.6,
  329.8,
  303.1,
  319.1,
  331.2,
  282.1,
  305.5,
  300.4,
  322.5,
  329,
  316.6,
  300.8,
  311.7,
  283.8,
  317.9,
  311.8,
  323.6,
  357.2,
  333.5,
  329.3,
  320.2,
  285.3,
  267.6,
  263.3,
  259.2,
  257.4,
  246.9,
  246.7,
  249.1,
  251.2,
  249.4,
  247.7,
  250.1,
  250.5,
  250.9,
  251,
  252.5,
  255.6,
  254.3,
  257.4,
  241.1,
  226.3,
  228.4,
  229.6,
  245.7,
  259.1,
  291.4,
  326.1,
  326.2,
  330.8,
  329.6,
  308.9,
  310.4,
  304.1,
  308,
  331.9,
  334.3,
  313.7,
  337.3,
  337.2,
  341.6,
  337.2,
  336.4,
  337.3,
  337.7,
  351.6,
  340,
  333.8,
  331.5,
  330.7,
  336,
  334,
  333.7,
  332.7,
  334.1,
  331.6,
  330.8,
  333.6,
  333.9,
  333.9,
  338.1,
  335.5,
  334,
  329.3,
  332.8,
  334.9,
  334,
  336.1,
  337.9,
  336.7,
  337.1,
  335.6,
  340.7,
  339.5,
  307.3,
  289.3,
  296.9,
  339.9,
  355.3,
  357.4,
  360.1,
  356.4,
  354.6,
  353.2,
  351.8,
  349.2,
  347,
  348.4,
  345.6,
  334,
  330.6,
  342.8,
  321.8,
  329.4,
  273.4,
  256.9,
  291.5,
  328,
  325.8,
  322.3,
  321.2,
  318.8,
  301,
  321.6,
  323.2,
  320.9,
  320,
  318,
  308.8,
  295.4,
  272.6,
  295.2,
  313,
  281.7,
  279.8,
  297.4,
  315.3,
  312.1,
  313.9,
  320.7,
  316.2,
  321,
  314.6,
  318.7,
  323,
  307.5,
  318.6,
  305.9,
  314.6,
  306.3,
  305.3,
  311.8,
  309.5,
  308.9,
  294,
  294.3,
  286.4,
  283.5,
  311.6,
  318.4,
  311.9,
  350.7,
  286.9,
  250,
  267.5,
  260,
  255.1,
  252.1,
  270.9,
  259.5,
  254.4,
  259,
  316.3,
  318.2,
  276.2,
  276,
  315.5,
  298.7,
  290.1,
  321.3,
  322.5,
  319,
  327.2,
  325.8,
  323.7,
  324.1,
  319.4,
  316.2,
  316.5,
  323.4,
  325.9,
  326.7,
  330.6,
  331.2,
  331,
  319.8,
  314.4,
  315,
  317.6,
  332.2,
  334.1,
  330.4,
  333.3,
  330.9,
  324.4,
  307.3,
  279.5,
  267.5,
  270.5,
  375,
  332.5,
  321.4,
  319.9,
  276.2,
  302.7,
  299.3,
  268.3,
  277.4,
  266.9,
  256.2,
  253.8,
  255,
  253.9,
  246.1,
  245,
  246.2,
  259.8,
  245.4,
  242.7,
  243.6,
  241.6,
  240.6,
  234.8,
  231.7,
  235.1,
  240.3,
  244.8,
  251.1,
  257,
  259.7,
  262.7,
  267.8,
  268.6,
  269.6,
  268.1,
  263.8,
  273.7,
  277.2,
  278.1,
  279.1,
  279.5,
  280.4,
  279.2,
  276.9,
  274.4,
  271.9,
  269.1,
  346.1,
  291.7,
  264.9,
  263.1,
  262.5,
  261.5,
  259.9,
  258.7,
  260.4,
  259.7,
  256.4,
  256.6,
  256.2,
  254.3,
  254.2,
  256.5,
  257.1,
  273.4,
  302.2,
  314.9,
  309.4,
  312,
  325.6,
  299.1,
  303.4,
  307.4,
  274.3,
  306.6,
  329.1,
  338.7,
  338.4,
  338.4,
  340.3,
  338.8,
  338.4,
  341,
  341,
  342.1,
  338.5,
  326.6,
  341.9,
  333.1,
  325.6,
  297,
  288.5,
  279.2,
  276.2,
  275.5,
  364.3,
  290.6,
  265.7,
  262.1,
  272.3,
  288.7,
  309.3,
  326.6,
  330.7,
  324.2,
  326.9,
  329.1,
  330.6,
  324.1,
  321.1,
  323.5,
  314.3,
  316.4,
  301.8,
  302.6,
  313.6,
  311.7,
  316.5,
  316.3,
  319.9,
  319.2,
  320.6,
  318.9,
  319.6,
  318.5,
  319.5,
  318.6,
  318.5,
  319.2,
  319,
  319,
  318.2,
  316.6,
  317.9,
  318.5,
  315.7,
  304.7,
  317.2,
  313.3,
  302.9,
  272.4,
  288.2,
  255.8,
  328.1,
  274.8,
  261.7,
  265.9,
  254.6,
  305.8,
  313.4,
  303.9,
  255.4,
  253.5,
  279,
  256.3,
  241.4,
  240.4,
  238.1,
  259.2,
  237.3,
  236.2,
  234.7,
  232.6,
  230.2,
  229.6,
  225.9,
  221.9,
  223.1,
  227.5,
  231.8,
  236.5,
  239.5,
  248.5,
  254.4,
  268.4,
  273.8,
  300.3,
  281.9,
  279.8,
  269.3,
  283.5,
  289.5,
  287.3,
  291.1,
  300.7,
  297.2,
  287.1,
  299.5,
  261.5,
  267.6,
  251.4,
  273.3,
  277.6,
  247.1,
  244.6,
  242.9,
  241.7,
  239.5,
  238.8,
  239.1,
  239.6,
  240.2,
  240.1,
  240.8,
  240.9,
  241.3,
  241.2,
  242.2,
  240,
  241.1,
  244.9,
  247,
  246.6,
  245.8,
  240.3,
  238.2,
  239.4,
  239.3,
  241.1,
  244.1,
  246.8,
  249.3,
  254.6,
  257.5,
  258.8,
  264.1,
  263.1,
  257.3,
  262.6,
  264.4,
  262.6,
  264.5,
  263.9,
  262.6,
  262.3,
  260.1,
  258,
  255.3,
  251.4,
  333.4,
  278,
  277.6,
  315.3,
  320.9,
  313.4,
  310,
  325.9,
  317.6,
  317.2,
  324.3,
  330.1,
  322.9,
  304.4,
  281.4,
  250.6,
  249.1,
  249.4,
  248.6,
  252,
  255.3,
  256.9,
  252.4,
  251.3,
  255.3,
  302.3,
  289.2,
  292.7,
  319.3,
  323.4,
  317.6,
  319.2,
  318.2,
  320.7,
  317.6,
  322.8,
  323.8,
  313.1,
  316.1,
  322.8,
  316.9,
  315.4,
  323.2,
  297.2,
  295.1,
  302.3,
  280.3,
  304.2,
  348,
  301.1,
  273.2,
  280.2,
  262.3,
  250,
  250,
  252.2,
  254.5,
  255.6,
  256.8,
  257.9,
  253.1,
  252.1,
  252,
  246.3,
  256.7,
  257.8,
  262.9,
  260.2,
  260.1,
  257.4,
  252.5,
  248.1,
  240.8,
  239.1,
  243.6,
  250.6,
  252.4,
  254.5,
  257.9,
  261.1,
  264.9,
  267.4,
  268.9,
  267.1,
  265.5,
  279.1,
  284.1,
  284.2,
  278.4,
  274.1,
  272.7,
  272,
  271.7,
  269.5,
  269.3,
  267.6,
  341.4,
  287.7,
  272,
  277.5,
  294.5,
  274.5,
  270.1,
  265.8,
  268,
  272.4,
  276.5,
  273.4,
  267.8,
  267.8,
  265.2,
  263.8,
  263.7,
  263.1,
  262.9,
  260.9,
  260.6,
  261.4,
  261.3,
  260.3,
  263.6,
  262.8,
  265.5,
  268.7,
  286,
  311,
  312.3,
  297,
  303.8,
  321.4,
  331.8,
  328.6,
  326.2,
  332.2,
  336.3,
  341.7,
  329.2,
  326.6,
  313,
  303.7,
  306.8,
  290.7,
  288.9,
  285.6,
  341.8,
  315.9,
  302.1,
  305.6,
  295.8,
  302.5,
  324.8,
  304.6,
  311.9,
  329.1,
  318.6,
  293.3,
  316.6,
  335.1,
  325.3,
  327.9,
  334.1,
  333.5,
  331.8,
  325.4,
  326.4,
  328.8,
  331.1,
  330.7,
  333,
  335.4,
  337,
  335.7,
  336.9,
  337.9,
  339,
  343.6,
  346.8,
  349.7,
  351.3,
  350.7,
  356,
  368.8,
  372.8,
  370.5,
  371.5,
  368,
  366.2,
  366,
  347,
  339.3,
  334.7,
  335.7,
  336.5,
  348.6,
  338.8,
  337.6,
  339.6,
  340.9,
  348.9,
  354.5,
  354.7,
  354.1,
  353.1,
  353.8,
  354.9,
  354.9,
  353.4,
  350.7,
  349.9,
  350.5,
  349.6,
  347.6,
  346.8,
  346.7,
  346.8,
  347.4,
  348.6,
  348.7,
  305,
  277.3,
  306.4,
  287.9,
  316.7,
  332.8,
  324.7,
  336,
  332,
  342.6,
  346,
  351.5,
  348.7,
  333.5,
  356.1,
  357,
  349.3,
  334.3,
  331.1,
  319.7,
  338.6,
  355.4,
  355.4,
  365.5,
  359,
  359.9,
  362.8,
  364.3,
  366.9,
  366.7,
  365.7,
  365.8,
  365.8,
  365.4,
  365.6,
  364.7,
  364.1,
  363.9,
  363.8,
  363.5,
  363.5,
  364,
  364.1,
  364.4,
  363.9,
  364.3,
  365.3,
  365.2,
  366.3,
  368.7,
  369.6,
  372.7,
  376.7,
  382.2,
  389,
  380.1,
  366.9,
  368.4,
  370.9,
  367.4,
  363.9,
  363.6,
  368.5,
  365.7,
  370.2,
  367.3,
  362.8,
  357.6,
  359.2,
  360.4,
  371,
  375.1,
  354.9,
  334.9,
  315.1,
  357.2,
  339.7,
  295.6,
  311.5,
  348.4,
  347.8,
  347.4,
  352,
  359,
  360,
  358.8,
  358.4,
  358.7,
  356.2,
  352.8,
  338.7,
  304.9,
  334.4,
  330.9,
  346,
  350.8,
  362.7,
  364.7,
  366,
  367.2,
  368.9,
  369.3,
  372.8,
  373.1,
  372.6,
  375,
  376,
  378,
  377.3,
  378.2,
  378.6,
  376.5,
  365.8,
  365.2,
  359.1,
  361.5,
  361.2,
  362.9,
  361.8,
  367.4,
  362.2,
  364.4,
  365.1,
  360.7,
  348.2,
  361.7,
  367.4,
  366.4,
  365.5,
  367.7,
  367.9,
  366.3,
  365.8,
  365.7,
  365.8,
  365.4,
  364,
  363.9,
  359.1,
  357.8,
  356.6,
  356.2,
  356.5,
  357.1,
  357.7,
  358.1,
  358,
  362.9,
  362.3,
  361.4,
  360.8,
  360.4,
  361.8,
  362,
  361,
  359.3,
  360.9,
  360.1,
  359.4,
  360.2,
  359.5,
  359.2,
  359.2,
  358.9,
  358.1,
  355.9,
  355.9,
  357.2,
  358.6,
  356.7,
  357.6,
  356.3,
  356.9,
  357.8,
  358,
  358.3,
  358.2,
  358,
  358.4,
  356.5,
  355.3,
  349.7,
  339.9,
  331.1,
  320.8,
  330.9,
  318.2,
  330.7,
  339.2,
  349,
  349.7,
  348.2,
  342.5,
  342.6,
  339.7,
  343.2,
  350.1,
  343.9,
  332.6,
  330.7,
  335.3,
  347.2,
  353.7,
  359,
  362.6,
  362.9,
  365,
  363.7,
  362.7,
  362.4,
  361,
  359.3,
  358.2,
  353.5,
  351.9,
  369.3,
  359,
  311,
  288.5,
  287.4,
  292.4,
  293.3,
  288.4,
  288.5,
  291.6,
  289,
  289.1,
  303.9,
  324,
  338.8,
  325.9,
  319.1,
  328.9,
  318.5,
  314,
  312,
  315.9,
  297.5,
  292.2,
  295.4,
  282,
  279.8,
  283.6,
  288.7,
  295.4,
  301.8,
  308.1,
  322.9,
  329.6,
  324,
  344,
  356,
  354.4,
  354.8,
  362.7,
  358.1,
  365,
  364.9,
  360.6,
  342.8,
  338.3,
  337.6,
  346.5,
  390.6,
  336.2,
  311.8,
  312.1,
  311.4,
  311.3,
  309.9,
  308.9,
  309.4,
  308.5,
  310.7,
  311.3,
  310.2,
  310.3,
  310.4,
  311.3,
  307.7,
  301.1,
  297.8,
  296.3,
  298.8,
  292.1,
  290.7,
  287.2,
  289.2,
  294.5,
  297.5,
  301.7,
  306.6,
  310.1,
  312.8,
  317.4,
  320.2,
  323,
  322.8,
  321.1,
  330.2,
  332.9,
  332.7,
  332.7,
  332.1,
  331.3,
  330.7,
  331.6,
  328.6,
  326.9,
  327.3,
  325.8,
  368.2,
  329.5,
  315.1,
  315.5,
  318.2,
  320.5,
  322.5,
  319.7,
  323.7,
  322,
  309.2,
  307.4,
  302.3,
  294.8,
  305.3,
  302.5,
  300.5,
  297.2,
  298.9,
  298.9,
  301.9,
  302.4,
  293.3,
  293.2,
  298.6,
  299.4,
  303.6,
  307.8,
  315.3,
  318.9,
  323,
  324.9,
  328.8,
  328.6,
  328.3,
  327.1,
  334.9,
  337.5,
  338.3,
  343.8,
  346.6,
  347.6,
  345.9,
  342.9,
  341.8,
  338.4,
  339.6,
  339.6,
  370.9,
  349.1,
  350.3,
  345.6,
  345.3,
  345.4,
  349.3,
  359,
  357.2,
  367.7,
  365.6,
  365,
  364.2,
  363.5,
  366.4,
  361.6,
  365.3,
  353.4,
  361.1,
  364.5,
  348,
  331.6,
  356.5,
  359.9,
  370.6,
  374.9,
  373.6,
  373.4,
  373.4,
  375.7,
  371.3,
  356.7,
  375.8,
  381.3,
  351.9,
  384.9,
  389,
  390.9,
  391.8,
  391.1,
  384.5,
  389.6,
  394.4,
  393.5,
  392.8,
  392.6,
  391.2,
  391.9,
  410,
  391.8,
  380.9,
  379.5,
  370.5,
  325.7,
  316.5,
  309.2,
  303.9,
  323.1,
  361.7,
  361.5,
  327.6,
  309.7,
  326.9,
  324.3,
  340.7,
  338.3,
  353.8,
  349.1,
  355.2,
  352.6,
  341.3,
  342.4,
  344.3,
  347,
  367.5,
  381,
  383.3,
  390.7,
  373.5,
  373.2,
  363.1,
  372.5,
  372.5,
  363.8,
  377.9,
  382.4,
  378.2,
  377.8,
  379.5,
  386.6,
  392.6,
  382.8,
  368.2,
  352,
  334.2,
  331.9,
  362,
  362.3,
  313.2,
  306,
  307.4,
  330.2,
  333.5,
  357.1,
  374.6,
  375.4,
  374.7,
  374.1,
  373.7,
  375.2,
  376.4,
  373.1,
  368.9,
  369.5,
  371.3,
  372.4,
  370.6,
  369,
  361.8,
  354.3,
  348.2,
  345.2,
  341.8,
  340.5,
  338.1,
  336.3,
  347.1,
  348.2,
  350.1,
  348.6,
  346.2,
  343.6,
  343.1,
  342.3,
  345.9,
  342.2,
  329.3,
  331.9,
  334.8,
  320.9,
  320.9,
  304.6,
  273.1,
  268.3,
  338.2,
  299.2,
  316.9,
  331.7,
  328.7,
  329.1,
  329.4,
  326.5,
  301,
  273.8,
  260.4,
  249.3,
  244.7,
  241.7,
  261.1,
  264,
  256.5,
  244.9,
  240.8,
  239.8,
  236.9,
  229.8,
  231,
  233.5,
  234.7,
  241.3,
  249.3,
  259.6,
  289.5,
  281.8,
  303.9,
  329.1,
  338,
  310.3,
  304.3,
  319.4,
  333.9,
  349.1,
  348.1,
  348.9,
  321.3,
  275.6,
  262.8,
  301.5,
  272.4,
  267.4,
  273.9,
  282.3,
  385.2,
  335,
  297.3,
  283.6,
  273.4,
  306.5,
  308.3,
  293.9,
  261.2,
  265.6,
  258.3,
  251.9,
  251.2,
  252.8,
  249.3,
  250.7,
  247.7,
  247.3,
  249.1,
  247.4,
  245.1,
  234.1,
  234.4,
  232.2,
  239.1,
  255,
  278.8,
  286,
  289.4,
  304.6,
  320.1,
  327.1,
  335.9,
  343,
  338.4,
  349.7,
  346.3,
  341.6,
  341,
  340,
  337.2,
  339,
  327.9,
  349.8,
  341,
  358.6,
  359.2,
  323.7,
  361.9,
  334.4,
  338.8,
  347,
  349.2,
  348.2,
  348.6,
  349.9,
  350.3,
  350.5,
  350.1,
  348.2,
  343.3,
  323.8,
  312.6,
  330.7,
  344.1,
  347,
  346.5,
  346.2,
  347.4,
  349.4,
  351,
  353.5,
  355.4,
  360.3,
  362,
  352.1,
  356.5,
  359.6,
  367.7,
  359.9,
  365.2,
  353.8,
  354.9,
  364.8,
  350.2,
  331.4,
  331.4,
  348.1,
  348.6,
  348.8,
  348.2,
  333.5,
  324.9,
  305.2,
  285,
  268.3,
  346.4,
  294.9,
  274.7,
  275.6,
  280.5,
  289.6,
  323.6,
  328.3,
  312.3,
  285.9,
  272.3,
  287,
  338.7,
  326.4,
  281,
  281,
  269.6,
  293.2,
  293,
  332.6,
  345.5,
  342.5,
  347.8,
  347,
  349.2,
  349.1,
  336.4,
  334.1,
  331.4,
  348.7,
  330.2,
  340.4,
  332.1,
  368.2,
  343.6,
  358.3,
  337.1,
  342.6,
  348,
  350.7,
  338.2,
  342.2,
  346.1,
  333.3,
  352.1,
  353.5,
  343.3,
  312.8,
  402.2,
  371.1,
  353.4,
  359.9,
  360.7,
  370.5,
  370.9,
  370.2,
  363.1,
  371,
  372.3,
  371.5,
  369,
  370.3,
  370.1,
  371.1,
  370.4,
  369.9,
  369,
  369.2,
  369.9,
  370.4,
  364.5,
  335.4,
  332.6,
  341,
  341.6,
  361.9,
  361.9,
  362,
  365.8,
  364.2,
  361,
  369.4,
  368.9,
  371.9,
  373.3,
  369.2,
  368.8,
  374.3,
  375.5,
  366.6,
  366,
  356.1,
  369.8,
  382,
  374.2,
  365.4,
  378.4,
  370.1,
  368.7,
  367.5,
  369,
  366.8,
  369.3,
  364,
  364,
  371.5,
  368.6,
  355.6,
  349.7,
  345.1,
  340.7,
  339.6,
  340.7,
  338.8,
  331.9,
  330.5,
  326.7,
  318.9,
  295.3,
  277,
  277.4,
  283.6,
  295.8,
  335,
  356,
  339.3,
  353.5,
  333.2,
  338.9,
  324.3,
  322.1,
  335.6,
  321.8,
  339,
  339.3,
  323.4,
  322.1,
  324.3,
  334.6,
  310.2,
  311,
  322.9,
  349.3,
  338.9,
  364.1,
  354.4,
  306,
  304.4,
  294.4,
  294.4,
  307.5,
  288.5,
  286.3,
  294.5,
  285.5,
  309.2,
  285.7,
  293.3,
  298.1,
  293.6,
  296.3,
  295.5,
  321,
  315.3,
  281.9,
  277.2,
  277.3,
  279.4,
  283.6,
  289.2,
  294.1,
  307.6,
  306.1,
  309.5,
  314.4,
  320,
  324.9,
  334.2,
  331.4,
  328.9,
  330.6,
  333.3,
  350.9,
  337.4,
  348,
  354.8,
  369.1,
  338.5,
  352.9,
  325.4,
  316.7,
  317.2,
  375.9,
  348.3,
  330.7,
  326,
  317.7,
  323.7,
  315.4,
  315.3,
  322.5,
  348.2,
  348.7,
  342.8,
  329.8,
  337.9,
  340.9,
  342,
  363.3,
  362.9,
  362.8,
  370.8,
  370,
  369.1,
  371.9,
  373.8,
  375.5,
  377.2,
  378.9,
  380.8,
  381.2,
  379.4,
  377.1,
  375.3,
  371.3,
  373.5,
  374.5,
  370.2,
  369.6,
  366.5,
  366.1,
  369.1,
  368,
  367.7,
  367.2,
  365.8,
  368.3,
  371.8,
  370.7,
  370.1,
  360.5,
  367.6,
  356.8,
  362.1,
  362.5,
  348.9,
  344,
  350.1,
  352.3,
  351.2,
  338.2,
  336.3,
  335.7,
  336.8,
  332.2,
  333.1,
  331,
  333.7,
  330.4,
  330,
  314.6,
  312.6,
  310.7,
  320.9,
  346.2,
  361.2,
  344.6,
  340.3,
  338,
  322,
  306.1,
  302.9,
  304.3,
  308.9,
  311.6,
  320.4,
  340.8,
  345.1,
  358.7,
  349.5,
  355,
  353.4,
  340.2,
  330.5,
  324.1,
  323,
  322.5,
  322,
  322,
  347.1,
  324.2,
  318.9,
  317.6,
  316.1,
  316.1,
  317.5,
  318.6,
  315.2,
  330.1,
  328.7,
  318,
  330.8,
  352.4,
  357.8,
  356.2,
  353.8,
  348.2,
  354.8,
  354.6,
  336.5,
  316.4,
  316.3,
  318.7,
  323.8,
  326.8,
  332.4,
  334.8,
  339.5,
  345.7,
  348.6,
  354.5,
  356.6,
  357.2,
  356.8,
  366.5,
  370.8,
  373.4,
  375.9,
  370,
  371.8,
  369.5,
  368.3,
  366.3,
  367.6,
  367.7,
  365.8,
  366.4,
  416.7,
  383.6,
  380,
  376.8,
  379.2,
  386.5,
  394,
  393.7,
  396.6,
  396.3,
  396.8,
  392.7,
  381.3,
  379.4,
  385.4,
  398.1,
  392,
  362.9,
  356.2,
  346.6,
  356.7,
  340.6,
  332.9,
  334.2,
  341.6,
  351.3,
  355.1,
  357,
  357.2,
  361.3,
  364.7,
  367.9,
  369.6,
  369.7,
  364.8,
  371.4,
  372.9,
  371.3,
  371.5,
  371.6,
  370.3,
  368.4,
  375,
  371.7,
  374.5,
  395,
  406.8,
  411.3,
  429.7,
  404.8,
  407.9,
  411.4,
  383.1,
  389.5,
  372.6,
  367.8,
  373.6,
  371.1,
  357.1,
  373.3,
  376.3,
  385.6,
  351.1,
  348.1,
  346.7,
  343.2,
  340.2,
  337.9,
  355.7,
  353.1,
  332.7,
  353.6,
  380.9,
  388,
  390.2,
  380.8,
  367.5,
  384.7,
  357.1,
  362,
  368.7,
  390.7,
  394.6,
  392.2,
  390.3,
  386.3,
  396.3,
  401.2,
  404,
  405.3,
  392.1,
  378.3,
  372.8,
  366.5,
  369.2,
  381.3,
  395.4,
  390.7,
  391.3,
  398.9,
  396.3,
  394.1,
  394.9,
  395.7,
  394.6,
  392.9,
  392,
  392.2,
  393.1,
  394.6,
  394.8,
  393.9,
  393.1,
  392.8,
  390.9,
  390.5,
  389.5,
  391.3,
  393,
  397.6,
  404,
  407.2,
  410,
  379.6,
  363.2,
  344.4,
  351.4,
  354.9,
  353.6,
  356.2,
  350,
  356.8,
  350.4,
  360.2,
  353.4,
  347.8,
  351.9,
  342,
  339.9,
  338.1,
  336.1,
  342.9,
  349.3,
  357.4,
  406.8,
  394.5,
  395,
  390,
  389.4,
  388.7,
  388,
  388.4,
  389,
  389.4,
  388.4,
  387.7,
  387.5,
  386.6,
  387.9,
  388.5,
  388.7,
  387.3,
  385.1,
  386.1,
  386.6,
  387.9,
  391.5,
  395.2,
  397.9,
  379.3,
  344.2,
  352,
  360.4,
  350.1,
  351.8,
  357.8,
  353.5,
  347,
  351.6,
  362.8,
  374.6,
  388.9,
  373.9,
  371.5,
  367.4,
  361.6,
  360.6,
  361.9,
  367.1,
  353,
  360.9,
  376,
  389.5,
  382.3,
  376,
  371.9,
  368.1,
  365.4,
  363.9,
  362.7,
  363.2,
  363.2,
  363.2,
  366.4,
  370,
  371.6,
  371.2,
  371.8,
  370.6,
  369.2,
  369.8,
  371.9,
  374.9,
  375.2,
  375.3,
  375.3,
  376.1,
  377.5,
  377.3,
  377.3,
  378.7,
  382.6,
  382.4,
  384.8,
  392,
  396.2,
  392.3,
  347.5,
  344.9,
  359.2,
  374.7,
  395.2,
  391.9,
  385.7,
  381.7,
  378.7,
  370.1,
  361.6,
  365,
  363.9,
  363.6,
  358.7,
  356,
  354.7,
  354.8,
  353.3,
  352.5,
  350.9,
  351.7,
  355.3,
  357.2,
  357.8,
  359.1,
  359.4,
  360.3,
  360.7,
  361.1,
  361.3,
  361.5,
  362.1,
  363,
  365.7,
  369.4,
  371.8,
  375.9,
  374.7,
  382.2,
  389.2,
  382.8,
  382.7,
  380.9,
  367.5,
  364.8,
  360.2,
  363.3,
  362.9,
  362,
  360.8,
  355.8,
  353.1,
  358.5,
  353.2,
  354.5,
  355.1,
  356,
  344.4,
  353.1,
  345.5,
  364.9,
  347.4,
  344,
  338.1,
  327.8,
  324.8,
  312.8,
  320.9,
  322.2,
  318.7,
  309.8,
  315.9,
  307.8,
  307.5,
  309.7,
  290.6,
  276.2,
  284.5,
  299.6,
  295.8,
  286.6,
  265,
  259,
  265.4,
  289.9,
  330.9,
  340.5,
  335.2,
  332.7,
  316.1,
  339.1,
  324.6,
  328.8,
  344.7,
  313.4,
  328,
  330.4,
  327.9,
  335.3,
  318.7,
  318.1,
  333.5,
  319.5,
  317,
  277,
  271.4,
  267.6,
  264.9,
  324.7,
  280.7,
  267.8,
  264.6,
  261.3,
  259.6,
  257.9,
  256.5,
  255.9,
  257,
  256.6,
  259.9,
  262.6,
  263.5,
  261.5,
  263.7,
  265.9,
  282.4,
  286.4,
  278.1,
  304.6,
  302.2,
  279.1,
  266.3,
  264.4,
  265.9,
  293,
  302.9,
  316.3,
  322.7,
  324,
  327.2,
  329.9,
  323.9,
  301.2,
  316.3,
  309,
  307,
  304.9,
  300.1,
  290,
  304.2,
  299.1,
  302.4,
  287,
  315,
  324.7,
  278.3,
  339.3,
  300.3,
  285.7,
  285.1,
  280.4,
  274.7,
  272.9,
  271,
  268.7,
  269,
  271.4,
  270.6,
  269.4,
  268.1,
  266.7,
  266.6,
  266.8,
  267.1,
  266.9,
  265.6,
  261.9,
  261.4,
  265.6,
  284.3,
  289.3,
  281.7,
  289.6,
  300.7,
  303.3,
  313.8,
  309.3,
  307.9,
  322.7,
  322.7,
  306.3,
  310.1,
  307.2,
  301.3,
  301.4,
  296.2,
  296.4,
  301.3,
  301.9,
  316.1,
  293.2,
  297.5,
  294.5,
  289.9,
  346.8,
  306.6,
  285.1,
  281.9,
  279,
  277.2,
  275.2,
  273.6,
  273.8,
  273.3,
  273.1,
  271.1,
  271.1,
  270.6,
  273,
  273.2,
  277.2,
  280.7,
  328,
  336.5,
  330.3,
  325.1,
  322.3,
  329.2,
  316.2,
  328.1,
  340,
  343,
  347.5,
  350.3,
  350.9,
  345.3,
  345,
  351.3,
  352.3,
  342.2,
  357.6,
  362.5,
  366.6,
  366.1,
  364.6,
  365.8,
  367.7,
  365.9,
  363.7,
  366.3,
  366.4,
  364.1,
  382.6,
  372.5,
  364.3,
  363.9,
  365.2,
  362.5,
  364.2,
  364.3,
  362.8,
  360.7,
  363.6,
  368.1,
  367.1,
  365.7,
  363.9,
  362.8,
  361.8,
  356.9,
  351.8,
  353.4,
  350.5,
  353.9,
  353,
  349.1,
  351.6,
  351.1,
  352.6,
  352.9,
  354.1,
  354.5,
  354.2,
  355.5,
  354.9,
  356.5,
  356.6,
  355.2,
  356,
  356.2,
  355.2,
  353.6,
  352.2,
  352.4,
  348.3,
  349.8,
  344.5,
  347.9,
  346.7,
  346.2,
  359,
  346.6,
  340.1,
  342.9,
  341.3,
  338.5,
  341.6,
  311.6,
  334.5,
  332.7,
  337.7,
  338.2,
  327.3,
  324.1,
  335.5,
  334.8,
  324.6,
  305.2,
  335.8,
  307.1,
  333.6,
  338.5,
  342.7,
  344.9,
  345.3,
  324.4,
  341.9,
  343.1,
  350,
  355.1,
  357.4,
  357.9,
  357.2,
  356.4,
  350.1,
  360.5,
  360.9,
  358.9,
  360.4,
  344.1,
  306.1,
  307.8,
  324,
  291.3,
  295.7,
  290.5,
  288.3,
  286.6,
  347.7,
  303.7,
  283.2,
  281.6,
  280.7,
  278.3,
  274.5,
  273.8,
  273.9,
  274.1,
  274.1,
  275.1,
  276.8,
  277.1,
  279.9,
  281.1,
  286,
  298.2,
  343.6,
  338.1,
  312.8,
  305.2,
  312.9,
  321.8,
  341.7,
  343.4,
  338,
  343.8,
  327,
  306.5,
  306.9,
  310.6,
  312.7,
  313.9,
  309.8,
  317.2,
  321.7,
  316.9,
  313.7,
  314.3,
  315.6,
  315.9,
  312.5,
  308.1,
  305.6,
  305.2,
  302,
  301.3,
  360.9,
  320.1,
  322.4,
  299.7,
  300.7,
  297.2,
  296.5,
  295.9,
  296.5,
  291.2,
  290.9,
  312.3,
  342.4,
  356.9,
  323.5,
  285.8,
  320.6,
  340.3,
  341.4,
  340.3,
  332.1,
  315.7,
  297.6,
  293.2,
  282.9,
  279,
  285.1,
  289.9,
  295.8,
  302.5,
  305.8,
  309.1,
  311,
  309.7,
  307.4,
  312.9,
  315,
  314.9,
  314.8,
  315.1,
  312.9,
  313.7,
  312.3,
  310.7,
  309.2,
  308.3,
  306.3,
  304.8,
  372.4,
  328.8,
  308.9,
  307.2,
  303.9,
  301.5,
  302.2,
  300.8,
  296.4,
  293.1,
  291.5,
  289,
  285.1,
  284.3,
  282.3,
  279.4,
  279,
  279.4,
  279.3,
  278.7,
  274.4,
  276.1,
  286.3,
  290.8,
  289,
  290,
  293.2,
  296.7,
  300.1,
  302.6,
  304,
  307.4,
  309.3,
  309.1,
  304.7,
  312.7,
  313.7,
  314.9,
  318.4,
  316.4,
  317.2,
  311.5,
  304.8,
  307.5,
  307.1,
  303.6,
  300.9,
  303.2,
  356.5,
  310,
  289.3,
  289.1,
  296.8,
  299.4,
  288.9,
  281.5,
  274,
  272.3,
  271.8,
  271.6,
  271.3,
  270.9,
  270.5,
  270.3,
  269.7,
  269.4,
  265.1,
  260.3,
  260.3,
  263.6,
  268.5,
  272.7,
  276.7,
  280.4,
  286.5,
  299.7,
  299.6,
  315.4,
  308.3,
  312.7,
  313.5,
  309.8,
  308,
  317.2,
  321.9,
  326.6,
  334.3,
  348.1,
  340.8,
  357.3,
  346.5,
  355.3,
  346.8,
  368.7,
  350.8,
  355,
  356.5,
  374.5,
  360.5,
  347.1,
  346.7,
  311.5,
  329.3,
  321.9,
  300.6,
  298.5,
  297.3,
  296.3,
  294.3,
  292.7,
  292,
  292.4,
  291.2,
  290.2,
  287,
  283,
  282.2,
  284.7,
  286.7,
  290.4,
  294,
  298.2,
  303.7,
  309,
  313.9,
  318.7,
  322.4,
  328.9,
  327.5,
  323.2,
  318.5,
  328.8,
  334.8,
  330.3,
  325.9,
  322.6,
  320.5,
  318.7,
  316.5,
  312.3,
  310.6,
  309.5,
  308.7,
  307.2,
  381,
  322.5,
  308.2,
  306.7,
  306.3,
  305.1,
  299.1,
  295.9,
  295,
  293.6,
  292.9,
  291.8,
  291.8,
  291.8,
  291,
  288.2,
  285.9,
  283.1,
  280.1,
  274.2,
  273.4,
  279.4,
  285.4,
  290.4,
  295,
  300.9,
  304.5,
  306.5,
  309,
  308.5,
  311.7,
  314.6,
  316,
  315.7,
  312.4,
  320.5,
  324.6,
  324.7,
  323.3,
  322.4,
  322,
  322.4,
  320.1,
  318.5,
  316.7,
  318.8,
  313.1,
  312.4,
  388.5,
  346.9,
  314.8,
  309.4,
  306.3,
  304.5,
  303.5,
  302.6,
  301.8,
  301.5,
  302.4,
  302.2,
  300.9,
  301.5,
  305.9,
  305.2,
  306.3,
  310.5,
  304.1,
  288.7,
  283.9,
  284.5,
  288.1,
  292.2,
  299.2,
  305.9,
  311.8,
  318.2,
  323.3,
  331.6,
  340.3,
  358,
  370.6,
  379.3,
  381.3,
  381.5,
  367,
  371.7,
  370.2,
  378.3,
  369.5,
  357.9,
  355,
  347,
  356.8,
  344.7,
  327.7,
  324.7,
  387.1,
  348.9,
  323.9,
  318.6,
  317.8,
  315.6,
  312.4,
  309.1,
  306.9,
  305.6,
  304.6,
  302.9,
  299.9,
  302.5,
  301.6,
  302.1,
  302.3,
  303.2,
  302.6,
  300.6,
  302.7,
  304.2,
  305.6,
  309.1,
  315.4,
  326.9,
  334.8,
  340.3,
  343.3,
  346.1,
  350.9,
  351.3,
  355.2,
  349.6,
  343,
  351.2,
  352.7,
  352.6,
  352.8,
  353.2,
  352,
  351.1,
  345.9,
  348.5,
  351.1,
  348.5,
  345.6,
  347.9,
  388.2,
  367.1,
  359.7,
  361.2,
  356.9,
  357.3,
  362.4,
  360.2,
  350.5,
  336.7,
  328.8,
  326.8,
  325.3,
  324.5,
  325.4,
  323.7,
  322.2,
  321.9,
  318.6,
  318.9,
  322.4,
  327.7,
  333,
  336.9,
  345.6,
  341.8,
  339.7,
  338.1,
  345.2,
  348.4,
  355.9,
  363.3,
  365.7,
  364.9,
  364.7,
  372,
  374.4,
  383,
  382.4,
  378.2,
  376.6,
  377.6,
  387.5,
  397.5,
  371.6,
  387.3,
  395.7,
  375.9,
  369.5,
  380.5,
  368.3,
  369.4,
  404.4,
  410,
  407.6,
  386,
  380.8,
  388.5,
  383.6,
  369.3,
  368.7,
  378.8,
  358.1,
  349.3,
  347.1,
  346.8,
  346.2,
  345.6,
  348.4,
  349.9,
  345.9,
  345.2,
  349.6,
  352.6,
  357.2,
  370.7,
  374.6,
  373.2,
  376,
  376,
  383.1,
  386.3,
  384.3,
  389.7,
  394.7,
  403.8,
  403.3,
  415.7,
  408.7,
  401,
  402.2,
  413.3,
  415.1,
  403.9,
  384.4,
  388.6,
  384.7,
  396,
  383.7,
  377.7,
  383,
  388.2,
  374.8,
  371.2,
  363.3,
  377.2,
  375.8,
  371.2,
  371.6,
  370.8,
  370.4,
  371.3,
  374.5,
  374.3,
  374.4,
  377.1,
  389.3,
  403.3,
  402.8,
  403,
  406,
  407.4,
  411.2,
  411.5,
  410.6,
  408.9,
  413,
  414.2,
  416.3,
  416,
  409.4,
  399.2,
  394.3,
  394.7,
  398.7,
  397.1,
  378.7,
  382.8,
  379.2,
  380.1,
  350.6,
  366.6,
  359,
  338.1,
  348.4,
  393.5,
  368.9,
  373,
  376,
  368.7,
  334.1,
  322.9,
  310.4,
  308.9,
  306.2,
  306.8,
  306.4,
  305.8,
  302.9,
  302.4,
  301.9,
  301.3,
  296.2,
  294.7,
  296.1,
  303.1,
  331.5,
  356.7,
  357.4,
  352.9,
  381.2,
  382.2,
  363.7,
  356.1,
  344.5,
  367.9,
  371.1,
  351.2,
  343.7,
  346.9,
  362.5,
  348.7,
  350.6,
  354.5,
  344.3,
  345.8,
  342.3,
  331.4,
  324.6,
  323.1,
  322.9,
  323.1,
  319.4,
  351.4,
  321.1,
  314.8,
  313.4,
  309,
  305.6,
  303.5,
  303.7,
  302.8,
  302.5,
  302.1,
  301.5,
  304.4,
  306.5,
  304,
  309.7,
  305.6,
  300.4,
  296,
  295,
  297.3,
  302.3,
  306,
  311,
  316,
  322.7,
  328,
  333.1,
  337.2,
  338.5,
  343.4,
  346,
  348.2,
  344.1,
  353.8,
  357.1,
  364.3,
  368,
  362.6,
  359.3,
  354.3,
  353,
  353.6,
  354.3,
  356.4,
  359.7,
  362.8,
  363.2,
  371.9,
  363.1,
  357,
  352.5,
  346.1,
  341.3,
  341.2,
  341.8,
  343.8,
  341.3,
  345.1,
  350.9,
  350.2,
  351.7,
  348,
  352.8,
  347.8,
  340.1,
  357.9,
  355.3,
  353.5,
  368.5,
  374.1,
  371.1,
  373.6,
  373.5,
  378.4,
  372.8,
  386,
  394.3,
  403,
  406.4,
  408.1,
  409,
  411.1,
  414.3,
  414.8,
  427.3,
  416.1,
  417.9,
  420,
  418.6,
  417.4,
  417.7,
  416.8,
  416.7,
  415.5,
  414.5,
  431.4,
  414.9,
  410.6,
  411,
  410.2,
  410.6,
  409.5,
  410.2,
  411.3,
  409.1,
  400,
  395.7,
  392,
  391.5,
  389.9,
  391.3,
  391.9,
  378.6,
  378.1,
  355,
  364.7,
  379.6,
  370.1,
  352.8,
  361.7,
  373,
  376,
  379.3,
  360.6,
  369.2,
  386.6,
  379.7,
  385.8,
  381,
  396.1,
  394.3,
  374,
  372,
  385.3,
  387.6,
  371.5,
  352.2,
  367.4,
  363.1,
  365.6,
  374.4,
  342.6,
  333.5,
  393.8,
  384.1,
  382.5,
  384.6,
  366.9,
  362.7,
  368.6,
  351.8,
  382,
  351.5,
  347.2,
  384.8,
  386.6,
  390.9,
  392.2,
  391.1,
  391.2,
  391.5,
  391,
  391.9,
  392.8,
  397.8,
  403.7,
  414.8,
  428.9,
  400.7,
  350.5,
  363.1,
  382.5,
  382.7,
  390.1,
  391.8,
  390.5,
  387.5,
  383.4,
  381.7,
  385.5,
  397.1,
  385.6,
  373.8,
  404.4,
  402.7,
  401.1,
  406,
  400.9,
  380.1,
  351.6,
  372.4,
  394,
  358.1,
  354.9,
  335.1,
  351.3,
  357.7,
  350.5,
  361.3,
  385.3,
  384.8,
  385.6,
  387.8,
  389.2,
  390.1,
  389,
  388.1,
  386.8,
  386.5,
  386.9,
  388.3,
  389.2,
  388.8,
  398.5,
  400.4,
  397.5,
  389.2,
  386,
  383.2,
  389.3,
  390.7,
  386.2,
  390.3,
  386.4,
  389.9,
  396.8,
  393.2,
  389.3,
  388.2,
  394.6,
  393.9,
  388.7,
  386.4,
  397.9,
  382,
  384.3,
  382.8,
  354.9,
  326.2,
  349.4,
  312.6,
  309.4,
  342,
  369.8,
  370,
  368.3,
  363.9,
  369.9,
  365,
  368.7,
  366,
  361.4,
  363.5,
  368.2,
  364.8,
  366.9,
  367.8,
  366.8,
  367,
  365.2,
  361.6,
  360.7,
  360.7,
  365.3,
  362.1,
  364.5,
  365.4,
  365.4,
  363.9,
  364.2,
  362.2,
  354.1,
  358,
  358.1,
  356.7,
  343.7,
  350.7,
  333.3,
  315.6,
  324.8,
  327.3,
  334.8,
  345,
  333.2,
  304.3,
  289,
  287.6,
  334.4,
  297.9,
  294.7,
  295.1,
  300.4,
  335.7,
  340.9,
  342.3,
  335.5,
  336,
  337.5,
  322.5,
  324.1,
  332,
  340.1,
  342,
  335.9,
  293.1,
  285.7,
  274.4,
  283.5,
  289.1,
  288.1,
  293.2,
  319.3,
  299.8,
  303.7,
  307.1,
  309,
  314.5,
  318.7,
  324.2,
  326.7,
  340.5,
  355.3,
  361.4,
  364.4,
  363.1,
  346,
  360.5,
  356.1,
  340,
  334.4,
  321.2,
  309.7,
  300,
  298.7,
  298,
  335.6,
  307.3,
  296.4,
  292.3,
  290.4,
  288.1,
  286,
  284.8,
  283.9,
  282.2,
  281.2,
  279.9,
  278,
  277.5,
  276.2,
  277.6,
  280.9,
  282.7,
  270.4,
  267.2,
  270.6,
  275.4,
  287.7,
  297.1,
  296.2,
  319.7,
  330,
  340.3,
  341.1,
  342,
  331.5,
  329.4,
  325.4,
  326.6,
  327,
  340.5,
  344.9,
  348,
  345.8,
  342.7,
  331.4,
  337,
  342.1,
  327.7,
  307.5,
  298.3,
  291.3,
  290.5,
  331.6,
  300.4,
  290.5,
  286.6,
  285.6,
  284.8,
  282.9,
  283.6,
  279.9,
  282.2,
  283.7,
  290.3,
  302.1,
  316.3,
  320.3,
  324.7,
  336.7,
  336.7,
  342,
  344.3,
  348.3,
  354.3,
  353.7,
  357.6,
  336.5,
  324.6,
  335.3,
  356.6,
  354.2,
  331.9,
  345.1,
  347.5,
  355.9,
  346.7,
  352.7,
  358.4,
  352.5,
  358.6,
  358.1,
  352.8,
  335.9,
  334.5,
  340.1,
  311.9,
  309,
  307.4,
  309.1,
  312.1,
  336.7,
  325.7,
  314.8,
  307.8,
  305.3,
  303.4,
  303.5,
  306.1,
  314.8,
  303.5,
  320.5,
  303.8,
  297.8,
  298.6,
  295.9,
  294.7,
  293.2,
  294.4,
  295.5,
  300.5,
  297.9,
  295.8,
  296.1,
  305.7,
  311.8,
  316.2,
  316.3,
  316,
  322,
  327.2,
  332.5,
  326.1,
  339.1,
  351.2,
  353.2,
  345.7,
  345.1,
  341.5,
  343.8,
  346.6,
  347.4,
  343.6,
  345.9,
  344.8,
  340.5,
  337.1,
  344.4,
  352.2,
  365.9,
  364.9,
  371.6,
  371.1,
  373.8,
  371.5,
  368.9,
  365.3,
  362.1,
  362.2,
  360.9,
  377.3,
  380,
  378.2,
  376.8,
  374.4,
  372.9,
  372.5,
  370.8,
  369.8,
  370,
  370,
  372.5,
  376.8,
  381.9,
  385.3,
  392.6,
  367.1,
  349.3,
  363.8,
  362.4,
  338.9,
  352.6,
  344.2,
  355.7,
  364.5,
  353.6,
  359.9,
  350.3,
  350.9,
  332.8,
  331.3,
  352.7,
  363.3,
  360.7,
  352.9,
  363.7,
  367.5,
  391,
  380.4,
  376,
  374.9,
  373.9,
  374.1,
  375.3,
  377.1,
  377.4,
  379,
  377.5,
  379,
  383.7,
  382.5,
  382.9,
  383.1,
  382.7,
  383.3,
  384.4,
  386.8,
  387.6,
  383.2,
  373.8,
  375.1,
  368,
  361.4,
  375.2,
  368.5,
  350.4,
  338.4,
  329.9,
  350.2,
  371.5,
  370.9,
  341.8,
  346.7,
  359.9,
  356.7,
  349.7,
  322.7,
  317.7,
  338.8,
  326.6,
  305.7,
  322,
  338.3,
  316.8,
  337.1,
  344.3,
  312.1,
  313.3,
  314.9,
  319.1,
  352.1,
  331.9,
  317.2,
  329,
  320.7,
  348.4,
  344.4,
  350.7,
  352.9,
  320.8,
  309.8,
  314.4,
  310.5,
  287.1,
  283.1,
  299.3,
  337.5,
  350.5,
  310.6,
  309.5,
  337.6,
  340.8,
  346.1,
  360.2,
  362.5,
  368.9,
  369.1,
  361.4,
  373.5,
  368,
  356.9,
  362.6,
  357.8,
  362.7,
  354.8,
  376.8,
  368.9,
  364.1,
  383,
  350.1,
  319.4,
  362.5,
  363,
  408.2,
  322.7,
  345.8,
  368,
  368.9,
  370,
  370.4,
  369.8,
  370.9,
  371.7,
  372,
  370.9,
  369.8,
  369.5,
  371.1,
  369.5,
  369.7,
  370.7,
  372.5,
  374.4,
  376.8,
  380.1,
  382.9,
  386.3,
  386.6,
  381.9,
  377.7,
  384.8,
  380.7,
  381,
  381.5,
  378.7,
  381,
  376.1,
  376.1,
  376.6,
  374.8,
  372.1,
  372.4,
  370.9,
  370.8,
  371.1,
  368,
  365.7,
  375.6,
  366.5,
  365.9,
  369,
  374.8,
  371.3,
  371.7,
  371.1,
  369.9,
  371.2,
  370.5,
  370.8,
  370.6,
  370,
  369.8,
  369.8,
  370.2,
  369.5,
  369.3,
  369.1,
  368.6,
  367.9,
  368.9,
  370.6,
  371.1,
  371.3,
  376,
  377.8,
  349.7,
  347.4,
  356,
  351.5,
  343.2,
  353.7,
  361.7,
  363.3,
  359.8,
  359.8,
  361.3,
  359.5,
  357.8,
  357.6,
  349.4,
  343.2,
  343.7,
  342.1,
  343.3,
  349.5,
  343.5,
  344.6,
  337.4,
  351.3,
  344.8,
  323.2,
  313.2,
  310.6,
  295.8,
  296.6,
  286.8,
  284.7,
  298.1,
  317.1,
  289.4,
  288.6,
  299.4,
  299.6,
  304.9,
  303.5,
  319.3,
  326,
  323,
  330.8,
  327.3,
  302.2,
  299.1,
  299.9,
  300.4,
  304,
  302,
  303.8,
  310.7,
  311.8,
  313.3,
  315.5,
  321.7,
  333.3,
  346.9,
  368.2,
  371.1,
  371.6,
  370.9,
  371.8,
  373.4,
  375.3,
  373.9,
  369.9,
  380.9,
  379.5,
  377.9,
  377,
  382.1,
  375.6,
  372.8,
  371.8,
  370.4,
  369.8,
  370,
  370.1,
  370.6,
  371.6,
  372,
  372,
  372.3,
  372.5,
  372.9,
  373.1,
  372.9,
  373.4,
  374,
  375.3,
  375.7,
  376.8,
  378.9,
  378,
  372.8,
  374.2,
  375.6,
  378.4,
  384,
  385.3,
  383.8,
  391.9,
  394.2,
  371.7,
  379.7,
  392.3,
  392.8,
  393.1,
  395,
  401.7,
  398.3,
  397.4,
  385.2,
  358.2,
  380.1,
  384.6,
  395.1,
  384.3,
  399.9,
  383.9,
  364.7,
  375,
  381.2,
  382.2,
  381.3,
  379.8,
  378.7,
  379.4,
  380.2,
  380.8,
  381.1,
  381.1,
  381.6,
  381.8,
  382.2,
  383.3,
  383.1,
  384.3,
  386.8,
  390.3,
  392.1,
  394.3,
  399.6,
  398.8,
  390.9,
  373.3,
  374.4,
  369.2,
  343.5,
  357.6,
  366.4,
  372.6,
  384.7,
  386,
  378.7,
  375.4,
  374.1,
  376.2,
  382.2,
  390.2,
  391.6,
  394.1,
  383.4,
  354.1,
  342,
  304.3,
  311.3,
  298.2,
  295.4,
  296.8,
  295.8,
  306.3,
  327,
  337.6,
  343.3,
  347.2,
  351,
  352.9,
  359.7,
  363.4,
  365.2,
  364,
  362.7,
  366.3,
  364.9,
  371.2,
  361.6,
  305.3,
  298.9,
  311.6,
  318.4,
  349.4,
  362.4,
  368.2,
  372.9,
  378.1,
  352.2,
  356.7,
  373.7,
  374.8,
  374,
  382.2,
  375.7,
  380.2,
  372.1,
  368.6,
  341.5,
  337.9,
  363.5,
  329.2,
  343.6,
  333.7,
  323,
  330.2,
  349.3,
  362.1,
  328.1,
  323,
  320.6,
  321.3,
  319.4,
  316.8,
  314,
  313.8,
  310.1,
  314.6,
  308.9,
  312.2,
  310.8,
  312.5,
  312.2,
  309.9,
  305.5,
  310.7,
  314.9,
  337.9,
  358.2,
  358.3,
  373,
  380.4,
  380.1,
  366.7,
  377.6,
  393.2,
  395.5,
  395.1,
  405.1,
  405.4,
  407.4,
  401,
  398.8,
  399.8,
  396.3,
  395.3,
  394.9,
  393.8,
  395.5,
  394.6,
  397.2,
  397.4,
  397,
  394,
  398.9,
  396,
  392.2,
  392.2,
  392.4,
  392.4,
  392.8,
  392.8,
  393,
  393.1,
  392.7,
  391.9,
  390.5,
  389.1,
  389,
  389,
  388.4,
  388.4,
  387.7,
  387.1,
  387.2,
  385.2,
  384,
  380.9,
  383.6,
  383.1,
  383.6,
  377.9,
  384.7,
  383.6,
  383.1,
  383.2,
  383.4,
  383.7,
  383.1,
  383.5,
  382.6,
  378.8,
  377.4,
  373.9,
  380.4,
  378.9,
  375.5,
  385.3,
  386.7,
  383,
  379.6,
  379.2,
  386.5,
  378.9,
  377.5,
  377.4,
  377,
  376.9,
  376.7,
  376.8,
  376.7,
  376.6,
  376.2,
  374.2,
  370.8,
  368.8,
  367,
  366.7,
  366.4,
  366.3,
  368.4,
  372.4,
  376.1,
  378.3,
  382.7,
  387.2,
  381,
  367.4,
  347.2,
  371.9,
  373.5,
  375.2,
  374.7,
  372.5,
  346.3,
  354.7,
  366.1,
  356.7,
  348.6,
  342.6,
  340.3,
  344.2,
  362.1,
  389,
  397.7,
  399.8,
  407,
  398.6,
  358.2,
  351,
  350.7,
  338.1,
  317.2,
  319.2,
  325.2,
  332.5,
  328.3,
  325.1,
  334.7,
  343.3,
  347.5,
  345,
  340.1,
  341.1,
  341.9,
  341.1,
  341.4,
  340.8,
  337.4,
  346.9,
  351.6,
  365.8,
  367.1,
  351,
  333.9,
  329,
  337.5,
  331.8,
  339.9,
  336.6,
  342.6,
  348.4,
  364.6,
  355.5,
  360.2,
  376.1,
  384.1,
  386.4,
  384,
  384.9,
  386.4,
  387.7,
  394.5,
  392.9,
  387.3,
  385.1,
  387.5,
  388.9,
  390.8,
  388.4,
  386,
  385.6,
  386,
  385.7,
  373.5,
  364.1,
  354.8,
  370.2,
  365.2,
  345,
  307.1,
  319.9,
  325.7,
  332.3,
  336.4,
  340.2,
  339.9,
  343.1,
  320.3,
  312.4,
  315.5,
  315.4,
  311.7,
  310.5,
  322.6,
  336.6,
  330.3,
  357.8,
  337.9,
  360.3,
  344.9,
  334.2,
  362.3,
  366.2,
  369.8,
  367.1,
  361.1,
  360.6,
  370,
  361.2,
  336.8,
  344.7,
  367.9,
  369.5,
  367.8,
  360,
  373,
  312,
  314.6,
  343,
  337.5,
  332,
  340.8,
  307.4,
  306,
  314.8,
  335.5,
  328,
  328.7,
  341.7,
  339,
  337.3,
  338.6,
  335.8,
  339.9,
  344.7,
  340.4,
  338,
  342.2,
  345.2,
  361.3,
  334.7,
  335.6,
  335.5,
  353.1,
  351.6,
  355.9,
  358.9,
  352.6,
  378.2,
  394.2,
  370.2,
  347.5,
  346.1,
  352.8,
  342.7,
  338.9,
  341,
  360,
  376.9,
  361.5,
  331.7,
  342.4,
  358.8,
  380.4,
  360.6,
  342.7,
  347.9,
  371.1,
  367.4,
  365.9,
  367.2,
  367,
  367.7,
  368.4,
  365,
  371.5,
  370.4,
  363.2,
  362.8,
  367.6,
  371.2,
  369.2,
  365.5,
  355.5,
  363,
  368,
  368.5,
  365.6,
  359.6,
  365.6,
  347.3,
  365.1,
  383,
  383.1,
  390.4,
  384.4,
  379.9,
  400.1,
  403.5,
  407.7,
  402.7,
  395.3,
  393.2,
  394.7,
  401.1,
  411.7,
  390.7,
  381.8,
  340.6,
  334.5,
  325.9,
  346.5,
  317.6,
  308.9,
  316,
  306.5,
  308.3,
  314.5,
  350.3,
  366.5,
  353.7,
  347.2,
  342.4,
  335.5,
  340,
  342.8,
  352.7,
  362.4,
  366.7,
  364.4,
  355.5,
  354.5,
  345.1,
  315.8,
  305.4,
  343.7,
  329.7,
  343,
  368.5,
  372.6,
  374.6,
  378.1,
  376.3,
  379,
  380.8,
  380.5,
  380.9,
  383.1,
  386.5,
  390.6,
  390.1,
  390.4,
  395.5,
  396.1,
  398.4,
  396.5,
  396.8,
  397.7,
  397.2,
  419.4,
  399.7,
  385.7,
  385.3,
  387.4,
  386.6,
  386.6,
  385.8,
  384.7,
  378.8,
  383.3,
  381.8,
  379.8,
  380.4,
  377.7,
  378.3,
  365.4,
  376.3,
  381.9,
  381.5,
  381.5,
  381.4,
  382.3,
  381.6,
  371.9,
  373.2,
  363.1,
  370.8,
  372.6,
  373.1,
  374.6,
  381.4,
  381.1,
  392.3,
  399.9,
  399.3,
  397.9,
  398.9,
  390.4,
  395.6,
  386,
  359.7,
  350.7,
  341.9,
  332.4,
  330,
  327.9,
  327.2,
  368.6,
  334.5,
  325.9,
  325.5,
  325,
  323.7,
  323.2,
  347.4,
  357.5,
  372,
  365.9,
  344.7,
  350.8,
  341,
  361.4,
  382.4,
  380.4,
  381.5,
  386.5,
  385.3,
  385.8,
  383.8,
  385.3,
  386.4,
  387.9,
  387.6,
  388.1,
  387.7,
  388.4,
  389.3,
  389.5,
  391.2,
  390.9,
  377.5,
  378.6,
  386.1,
  392.9,
  387.4,
  382.8,
  378.1,
  376.7,
  382.7,
  375.7,
  362.4,
  357.1,
  350.5,
  348.5,
  336.8,
  370.8,
  337.3,
  330.4,
  328.5,
  324.4,
  320.8,
  318,
  322.5,
  370.9,
  380.8,
  382.3,
  382.9,
  383.9,
  384.1,
  383.5,
  382.3,
  381.9,
  381.8,
  382.1,
  381.4,
  380.9,
  381.2,
  381.2,
  381.5,
  383.2,
  384.8,
  385.7,
  387.4,
  388.2,
  388.4,
  388.5,
  389.2,
  386.1,
  391.6,
  393,
  394.8,
  395.2,
  386.1,
  382.2,
  376.1,
  356.1,
  362.2,
  353.3,
  354.1,
  352.1,
  335.5,
  323.4,
  320.1,
  370.1,
  328.9,
  314.8,
  311.7,
  308.7,
  305.9,
  304.5,
  304.8,
  311.3,
  325.3,
  335.5,
  341.8,
  346.6,
  349.1,
  359.2,
  362,
  363.5,
  368.9,
  373.4,
  378.2,
  382,
  384.5,
  386.7,
  388.9,
  389.1,
  381.4,
  333.1,
  329.2,
  336.6,
  340.1,
  345.1,
  360,
  369.6,
  371.5,
  366.9,
  371.5,
  374.2,
  383.2,
  393,
  378.5,
  387.6,
  356.9,
  365.4,
  348.1,
  361.5,
  344.6,
  341,
  341.2,
  364,
  346.2,
  337,
  332.7,
  331.8,
  331.1,
  328.6,
  326.7,
  325.3,
  324.5,
  323.1,
  322.4,
  322.8,
  321.1,
  321.2,
  321.6,
  322.4,
  320.3,
  319.4,
  322.7,
  316.4,
  318.5,
  322,
  327.9,
  332.4,
  338.5,
  342.8,
  347.1,
  349.4,
  350.6,
  354.6,
  360.8,
  370.1,
  371.9,
  370.6,
  383.9,
  386.2,
  383.7,
  378.6,
  390.8,
  370.8,
  385.9,
  379.1,
  354.3,
  350.8,
  349.3,
  348.7,
  348.5,
  376.5,
  352.9,
  348.9,
  347.9,
  342.1,
  347.8,
  372.2,
  364.8,
  338.8,
  340.4,
  358.3,
  348.5,
  358.8,
  346.6,
  367.2,
  369.9,
  389.5,
  389,
  385.4,
  383.1,
  386.9,
  386.6,
  388.8,
  388.5,
  387.1,
  391.5,
  393.9,
  387.7,
  372,
  367.7,
  370.1,
  366.9,
  372,
  375.4,
  384.5,
  388,
  402.5,
  414.1,
  411.5,
  411.7,
  404.4,
  376,
  363.8,
  359.9,
  357.6,
  353,
  351.4,
  350.1,
  378.2,
  351.4,
  345.2,
  377.9,
  383.9,
  387.2,
  382.9,
  363.8,
  340.7,
  341.9,
  352.1,
  362.3,
  370,
  378.2,
  380.9,
  383.8,
  383.6,
  384.8,
  384.1,
  383.6,
  386.6,
  395.8,
  405.9,
  387.1,
  346,
  366.2,
  378.9,
  382.6,
  365.7,
  381.8,
  398.4,
  400.2,
  385.8,
  376,
  385.8,
  395.9,
  388.2,
  383.9,
  374.6,
  379.6,
  376.1,
  398.8,
  404.3,
  397.2,
  397,
  407.2,
  404.2,
  387.9,
  421.7,
  395.9,
  376.8,
  371.1,
  379.6,
  387.3,
  386.4,
  388.4,
  388,
  392.2,
  388.4,
  383.1,
  383.4,
  383.6,
  384.4,
  381.3,
  382.6,
  391,
  385.8,
  383.4,
  386.9,
  391.4,
  384.4,
  377.4,
  351.1,
  352.5,
  355.6,
  384.6,
  375.9,
  364.8,
  361.5,
  357.1,
  355.7,
  355,
  391.7,
  386.5,
  390.8,
  393.2,
  399.2,
  387.2,
  382.7,
  368.8,
  374.8,
  366.7,
  364.5,
  337.7,
  330.9,
  328.7,
  342,
  329.4,
  330.9,
  332.6,
  333.7,
  327.4,
  328.3,
  335.7,
  344.2,
  359.4,
  371.1,
  372.5,
  375.2,
  368.7,
  360.5,
  361.1,
  365.6,
  371.6,
  372.1,
  383.1,
  383.2,
  385.4,
  380.9,
  386.5,
  394.2,
  379.1,
  362.2,
  381.8,
  378.9,
  393.5,
  393.4,
  388.5,
  382,
  382.9,
  384.1,
  380.8,
  374.6,
  358.8,
  359.7,
  369,
  394.9,
  390.3,
  396.3,
  400,
  403.2,
  403.9,
  367.6,
  343.6,
  364.5,
  347.5,
  354,
  354.7,
  345.9,
  341.1,
  340.7,
  338.1,
  338.6,
  360.2,
  365.6,
  369.8,
  376.6,
  382,
  383.1,
  384.6,
  389.5,
  389.2,
  389.1,
  389.7,
  391.9,
  395.7,
  401.2,
  408.2,
  411.1,
  408.5,
  407.6,
  406.1,
  408.2,
  418.9,
  426,
  415.5,
  398.1,
  393.1,
  389.2,
  392.9,
  379.6,
  382.3,
  373,
  375,
  384.3,
  378.2,
  379.9,
  381.8,
  378.3,
  349.2,
  372.4,
  404.7,
  394.1,
  384.8,
  382.3,
  384.6,
  383.5,
  381.7,
  381.9,
  380.7,
  381.1,
  381.2,
  381.2,
  381,
  380.9,
  384.6,
  381.1,
  378.5,
  377.3,
  381.9,
  371.9,
  372.1,
  372.8,
  360.4,
  337.4,
  348.2,
  344.6,
  355.7,
  372.9,
  379.8,
  376.4,
  376.2,
  383.6,
  384,
  372.4,
  384.6,
  392.3,
  391.3,
  390.5,
  402.7,
  389.5,
  385.2,
  382.2,
  389.6,
  395.5,
  394.4,
  393.9,
  393.5,
  393.1,
  401.1,
  395.4,
  389.3,
  387.9,
  386.3,
  383.7,
  383.1,
  382.9,
  382.4,
  381.8,
  381.1,
  380.3,
  382,
  382.4,
  382.2,
  381.4,
  381.1,
  380.9,
  380,
  379.9,
  380.1,
  382,
  386.1,
  392.8,
  397.6,
  399.2,
  399.6,
  405.8,
  415.4,
  421.5,
  431.4,
  409.6,
  370.4,
  388.5,
  386.1,
  408.2,
  409.5,
  407.4,
  408.4,
  396.7,
  406.3,
  408.5,
  410.9,
  413.7,
  408.6,
  409,
  404.9,
  401.7,
  425.1,
  413.4,
  404.1,
  395.1,
  391.5,
  382.4,
  379.6,
  379.2,
  378.1,
  378.2,
  378.2,
  378.7,
  378.5,
  379.7,
  380.3,
  379.4,
  379.7,
  379.4,
  379.7,
  378.3,
  379.9,
  384.1,
  392.4,
  395.3,
  397.6,
  373.8,
  329.9,
  335.6,
  338.3,
  346.6,
  359.1,
  365.7,
  371.4,
  369.3,
  384.9,
  386.1,
  389.3,
  382.9,
  377.1,
  371.9,
  369.3,
  351.4,
  336.4,
  331.8,
  329.1,
  342.3,
  324.9,
  327,
  439,
  421.2,
  366.9,
  336.2,
  329,
  331.1,
  344.5,
  351.6,
  368.8,
  375.6,
  374.4,
  368.5,
  365,
  370.1,
  377.4,
  378.7,
  377.9,
  377.3,
  377.5,
  377.4,
  376.9,
  380,
  383.6,
  386.5,
  374.3,
  346.7,
  350.5,
  366.7,
  359.4,
  349,
  360.5,
  362.4,
  352.1,
  376.4,
  390.5,
  376,
  390.8,
  395.2,
  379.5,
  402.7,
  402.3,
  404.7,
  407.3,
  398.1,
  397.8,
  380.4,
  340.4,
  336.2,
  415.5,
  360.4,
  342.1,
  340.1,
  344.2,
  335.5,
  345.6,
  362.5,
  365.4,
  365.7,
  369.5,
  358.6,
  349.3,
  364.5,
  365.7,
  360,
  352.2,
  351.6,
  365,
  373.5,
  373.3,
  374.2,
  378,
  379.3,
  376,
  371.6,
  369,
  381.5,
  379.4,
  380.6,
  382.9,
  387.8,
  395.3,
  395.2,
  396.9,
  399.1,
  402,
  409.7,
  405.9,
  405.6,
  410.6,
  407.2,
  409,
  408.6,
  406.6,
  407,
  404.3,
  402.7,
  409.4,
  402.5,
  402,
  402.5,
  402.6,
  402.5,
  403.8,
  403.7,
  403.5,
  404,
  404.6,
  405,
  404.4,
  404.5,
  403.2,
  400.4,
  398.6,
  397.6,
  397.3,
  396.7,
  398.2,
  398.1,
  400.9,
  402.7,
  408.4,
  409.7,
  408.1,
  398.2,
  402.7,
  400.5,
  401.9,
  385.5,
  384.2,
  388.3,
  389.2,
  404.2,
  410.1,
  406.5,
  399.9,
  399.9,
  395.7,
  409.2,
  401,
  370.1,
  353.3,
  352.9,
  361.5,
  354.3,
  392.4,
  360.2,
  339.5,
  339,
  335,
  333.4,
  335.7,
  346.3,
  355.6,
  363,
  368,
  369.6,
  374.4,
  374.9,
  384.4,
  388.7,
  389.3,
  387.1,
  379.7,
  372.4,
  365.4,
  357.6,
  361.8,
  359.3,
  316.2,
  320.7,
  342.8,
  340.2,
  346.4,
  339,
  347.6,
  356.2,
  368.8,
  369.8,
  366.3,
  362.1,
  364.7,
  355.2,
  350.8,
  355.9,
  349.7,
  342.5,
  340.1,
  338.1,
  335.7,
  336.2,
  335.6,
  336.6,
  378.8,
  366.6,
  338.1,
  341.4,
  345.2,
  352.7,
  338.2,
  333.1,
  337.6,
  338.2,
  332.9,
  330.4,
  332.7,
  341.2,
  334.9,
  331.4,
  331,
  339.7,
  331.9,
  326.7,
  321.5,
  313.6,
  319.7,
  332.9,
  355.4,
  367.2,
  369.7,
  376.7,
  381.9,
  385.7,
  386.2,
  388.5,
  389.3,
  392.1,
  400.3,
  393.1,
  403.6,
  408.1,
  411.6,
  413.5,
  417.7,
  419.6,
  399.1,
  365.6,
  361.4,
  368.1,
  370.8,
  379.9,
  413.3,
  395.7,
  389,
  389.7,
  383.6,
  360.1,
  347.8,
  338.3,
  331.5,
  363,
  375,
  379.5,
  376.8,
  379,
  387.6,
  381.1,
  381.6,
  374.1,
  371.2,
  382.1,
  390.1,
  390.7,
  390.7,
  390.3,
  392.2,
  397.1,
  397.3,
  394.1,
  390.1,
  391.1,
  400.6,
  384.2,
  392.5,
  388.6,
  377.3,
  394.1,
  387,
  381.4,
  386.2,
  385,
  378.2,
  386.5,
  388.1,
  388.3,
  384.2,
  375.4,
  362.6,
  370.2,
  379.2,
  368.8,
  343.7,
  324.8,
  329.5,
  316.8,
  326.3,
  338.2,
  372.6,
  379.1,
  381.4,
  380.9,
  380.9,
  381.3,
  382.6,
  384.1,
  383,
  381.9,
  384.3,
  381.4,
  333.3,
  358.9,
  319.2,
  343,
  348,
  328.2,
  352.4,
  334.2,
  343.5,
  348.8,
  365.2,
  359.9,
  362.9,
  359.8,
  368,
  361.9,
  379.9,
  373.9,
  359.6,
  363.5,
  371,
  380.7,
  386.4,
  380,
  385.5,
  395,
  398.7,
  397.9,
  400.5,
  399.2,
  398.4,
  395.8,
  397.1,
  401,
  399.5,
  399.2,
  399.6,
  400.5,
  400.7,
  401.5,
  403.5,
  404.5,
  405.2,
  402.1,
  400.3,
  400.2,
  398.6,
  399,
  400,
  399.6,
  399.5,
  400.5,
  400.4,
  397.5,
  398,
  379.1,
  391.1,
  389.5,
  387.5,
  387.6,
  383.8,
  386.6,
  386.7,
  385.5,
  384,
  385.4,
  374,
  356.8,
  355.4,
  369.9,
  365.3,
  367.4,
  344.7,
  341.1,
  327.4,
  313.5,
  367.8,
  328.9,
  317.1,
  312.3,
  313.5,
  311,
  312.8,
  327.5,
  335.6,
  341.8,
  342.7,
  347.9,
  353.1,
  355.9,
  350.8,
  348.7,
  346.2,
  345.6,
  345.8,
  346.8,
  349.3,
  342,
  331.9,
  341.2,
  354.9,
  331.2,
  323.9,
  330,
  333.8,
  339.3,
  356.9,
  354.5,
  355.1,
  377.8,
  372.7,
  368.6,
  371.9,
  368.5,
  384.2,
  391.2,
  387.1,
  386.1,
  380.4,
  374,
  358.1,
  340.4,
  336.4,
  331.8,
  371.6,
  343.7,
  341.7,
  333.5,
  333,
  331,
  330.7,
  330.9,
  333.5,
  338.3,
  347.4,
  345.1,
  343.4,
  350.2,
  354.3,
  357.6,
  360.3,
  359.1,
  353.5,
  349.3,
  346.2,
  347.4,
  345.4,
  322.6,
  315.2,
  320.3,
  326.3,
  331.9,
  338.4,
  344.3,
  348.4,
  355.7,
  359.9,
  365.8,
  366.2,
  368.6,
  362.7,
  364.8,
  362.7,
  363.9,
  359,
  363.3,
  362.6,
  357,
  350.4,
  349.1,
  349.1,
  352.4,
  379,
  364.5,
  355.8,
  349.1,
  347.8,
  343.5,
  339.8,
  337.3,
  337.9,
  332.5,
  327.8,
  328.1,
  326,
  328.3,
  328.1,
  327.4,
  327.4,
  329.2,
  329,
  327.4,
  331.3,
  324.6,
  325.2,
  325.6,
  333.3,
  348.1,
  367.5,
  369.5,
  381.8,
  366.8,
  373.6,
  396,
  401.3,
  402.6,
  406.1,
  408.3,
  420.2,
  406.6,
  405.2,
  404.3,
  401.5,
  396.8,
  396,
  373.4,
  378.5,
  382.4,
  339,
  326,
  370,
  323.2,
  318,
  318.3,
  337,
  335.8,
  344,
  334.6,
  336.4,
  348.9,
  350.8,
  347.8,
  347.8,
  352.2,
  355.8,
  358.2,
  360.9,
  359.3,
  364.8,
  359.7,
  352.2,
  361.5,
  372.6,
  356.9,
  340.2,
  334.6,
  367.1,
  378.8,
  385.4,
  379.4,
  371.4,
  374.1,
  368.2,
  363.8,
  372.8,
  370,
  372.6,
  375.8,
  383.2,
  378.5,
  374.7,
  369.7,
  377.7,
  374.5,
  373,
  374.2,
  365.5,
  370.7,
  384,
  371.6,
  367,
  373.8,
  376.5,
  383.3,
  383.5,
  383.3,
  383.3,
  383.5,
  383.5,
  384.3,
  384.3,
  384.3,
  384.3,
  385.2,
  385.4,
  385.4,
  385.2,
  385.3,
  385.5,
  386.2,
  387.1,
  388.7,
  390.5,
  394.5,
  397.4,
  399.3,
  401.3,
  413,
  425,
  425,
  382.5,
  389.8,
  378.9,
  390.1,
  389.7,
  385.4,
  390,
  387.3,
  386.3,
  389.5,
  392.7,
  394.1,
  389.7,
  387.6,
  389.4,
  392.5,
  395.3,
  401.5,
  399.3,
  397.8,
  397.8,
  398,
  397.3,
  396.8,
  397.1,
  397.2,
  398.1,
  398,
  398.5,
  399.1,
  399.6,
  400.1,
  400.8,
  401.4,
  401.4,
  401.9,
  403.2,
  403.9,
  405.9,
  408.7,
  409.3,
  412.1,
  417,
  423.4,
  441,
  398.5,
  372.6,
  380.1,
  378.2,
  389.5,
  376.8,
  380.2,
  372.9,
  379,
  367.5,
  370.2,
  381.2,
  373.3,
  358.5,
  349.2,
  342.1,
  337.6,
  334.4,
  353.6,
  388.5,
  350.3,
  340.1,
  338.4,
  333.4,
  332,
  333.3,
  328,
  331.4,
  358.2,
  335.2,
  340.3,
  338.6,
  334.2,
  327.9,
  334.6,
  348.4,
  374.6,
  372.9,
  363.3,
  345.3,
  334.2,
  336.7,
  335.7,
  343.7,
  350,
  332.3,
  350.1,
  350.8,
  364,
  372.1,
  386.3,
  386.8,
  382.6,
  366.7,
  377.7,
  390.2,
  392.8,
  397.1,
  400,
  400.2,
  399.9,
  399.9,
  399.9,
  399.8,
  400,
  399.9,
  398.7,
  405.9,
  393.8,
  390.4,
  363.2,
  362.7,
  377.6,
  379.4,
  366.6,
  362.8,
  353.3,
  344,
  349.3,
  369.8,
  334.7,
  326.5,
  327.7,
  354,
  359,
  352.5,
  366.7,
  362,
  334.2,
  327.5,
  338.4,
  373.7,
  364.2,
  339.8,
  338.1,
  338.2,
  346.8,
  354.3,
  347.4,
  349,
  348.2,
  345.1,
  359.2,
  378,
  391.9,
  396.5,
  406.6,
  403.9,
  398.2,
  389.6,
  373.1,
  361.7,
  338.2,
  333.3,
  332.5,
  360.9,
  331.8,
  322.8,
  319.4,
  316.3,
  314.3,
  312.3,
  310.6,
  309.5,
  308.4,
  306.4,
  305.1,
  303.9,
  302.1,
  299.4,
  297.6,
  298.6,
  299.2,
  294.8,
  294.8,
  291.4,
  294.9,
  300.7,
  306,
  315.3,
  317.5,
  321.8,
  321.3,
  320.2,
  321.6,
  321.7,
  328.9,
  330.1,
  333.2,
  327.9,
  337.4,
  344,
  348.8,
  356.5,
  355.4,
  346.7,
  348.9,
  350.3,
  341.5,
  340.1,
  342.5,
  345.1,
  334.9,
  372,
  340,
  337.3,
  335.9,
  333.8,
  328.6,
  325.1,
  323.3,
  322.1,
  319.9,
  318.7,
  319.8,
  322.2,
  324.8,
  324.9,
  324.8,
  324.4,
  323.3,
  322.5,
  321.1,
  315.3,
  314.1,
  316.9,
  320,
  324.4,
  329.9,
  335.5,
  340.2,
  347,
  352.1,
  356.1,
  358.2,
  357.1,
  356.1,
  354.1,
  365.7,
  366.4,
  372.6,
  374.3,
  369,
  365.6,
  366.1,
  360.5,
  356.2,
  355.1,
  353.8,
  352,
  432.5,
  380.9,
  351.8,
  347.4,
  346.7,
  345.3,
  344.9,
  345.2,
  343.8,
  342.3,
  341.6,
  340.9,
  338.7,
  336,
  334.6,
  333.5,
  330.3,
  329.4,
  328.1,
  327.1,
  326.4,
  323.2,
  322.2,
  325.7,
  328.3,
  332,
  337.9,
  342.8,
  346.3,
  349.2,
  351.5,
  357,
  360.4,
  362.4,
  365.1,
  356.7,
  366.2,
  375.3,
  378.9,
  378,
  381.8,
  378,
  379.5,
  372.5,
  374.7,
  370.1,
  363.6,
  361.5,
  433.9,
  384.5,
  356.9,
  353.2,
  354,
  354.2,
  354.6,
  353,
  352.4,
  350.2,
  346.3,
  345.3,
  345.9,
  353.1,
  361.8,
  360,
  347.9,
  343.7,
  349.2,
  340.2,
  336.2,
  334.1,
  329,
  330.2,
  332.4,
  335.6,
  340.9,
  347.4,
  353.6,
  356.2,
  362.2,
  365.1,
  368.3,
  369.3,
  368.5,
  362.7,
  372.5,
  379.6,
  387.3,
  392.9,
  380.2,
  387.8,
  385.6,
  384.6,
  377.3,
  367,
  366.5,
  366.3,
  425.1,
  386.3,
  369.1,
  366.1,
  364.5,
  366.7,
  365.1,
  362.2,
  361.2,
  357.7,
  358.7,
  355.5,
  353.1,
  353.6,
  353.8,
  355.5,
  354.4,
  350.4,
  348,
  346.1,
  345.6,
  340.3,
  333.8,
  334.3,
  337.7,
  342,
  348.3,
  356.2,
  359.9,
  366.9,
  371.8,
  378,
  386.1,
  393.3,
  399.6,
  410.9,
  407.6,
  401.2,
  400.2,
  400,
  412.8,
  418.4,
  423.5,
  422,
  411.6,
  401,
  386.9,
  383.6,
  425.6,
  400.8,
  374.8,
  374.3,
  368.5,
  370.5,
  369,
  363.7,
  365.2,
  369.8,
  364,
  366.7,
  368.6,
  370.7,
  365.5,
  372,
  382.4,
  384.3,
  379.4,
  376.3,
  375.8,
  365.7,
  360.2,
  352.5,
  344.2,
  348.3,
  353.2,
  359.1,
  363.7,
  368.5,
  374.6,
  379.6,
  384.4,
  385,
  390,
  389.3,
  391,
  387.8,
  389.1,
  389.6,
  392.1,
  381.1,
  377.7,
  377.8,
  375.7,
  375.2,
  377.1,
  377.1,
  437.1,
  399.2,
  373.1,
  385.1,
  379.7,
  378.5,
  369.5,
  363.5,
  358.3,
  355.8,
  357.5,
  357.4,
  354.5,
  353.3,
  352.2,
  349.6,
  348.3,
  348.4,
  346.2,
  345.1,
  343.9,
  334.5,
  329,
  327.9,
  329.8,
  331.6,
  334.2,
  342.1,
  352,
  356.7,
  359.1,
  360.7,
  363.7,
  367.3,
  369,
  362.1,
  370.6,
  374.8,
  375.8,
  376,
  375.7,
  373.1,
  371.8,
  369.9,
  367.4,
  365.7,
  366.4,
  364.4,
  428.2,
  382.7,
  364.5,
  362.6,
  362,
  361.6,
  358.6,
  355.3,
  353.4,
  351.7,
  351,
  350.2,
  350.8,
  351.1,
  349.8,
  349.1,
  347.3,
  346.4,
  346.4,
  345,
  342.7,
  335.5,
  331.2,
  332.3,
  335.7,
  339.9,
  346.6,
  351.5,
  356.1,
  361.3,
  366.1,
  372,
  376.6,
  378.1,
  375.1,
  370.9,
  377.2,
  382.3,
  381.7,
  378.5,
  378.7,
  377.9,
  376.4,
  378.9,
  380.1,
  378.7,
  377.9,
  375.5,
  445.2,
  401.8,
  374.2,
  373,
  373.4,
  375.3,
  374.8,
  372.2,
  371.4,
  368.2,
  365.5,
  361.2,
  363.6,
  364.4,
  364.1,
  365.3,
  360.9,
  358.5,
  356.1,
  359.2,
  357.9,
  355.4,
  347.4,
  341.2,
  344.2,
  348.5,
  354.3,
  359.8,
  365.1,
  370.4,
  376.3,
  377.9,
  380.6,
  381.3,
  380.1,
  375.4,
  382.1,
  386.1,
  384.7,
  388,
  386.7,
  388.2,
  392,
  397,
  396.8,
  395.5,
  397.3,
  403.4,
  435.3,
  413,
  386.7,
  377.3,
  371.1,
  362.5,
  359.2,
  355.2,
  352.6,
  350.6,
  350.5,
  350.5,
  348,
  344.3,
  341.2,
  340,
  338.4,
  338.5,
  337.3,
  334.9,
  334.8,
  337.7,
  386.1,
  393.2,
  398.1,
  399.1,
  399.7,
  400.8,
  402.6,
  398,
  391.9,
  407.6,
  409.5,
  411.2,
  411.1,
  411.2,
  412.7,
  413.2,
  410.4,
  410,
  408.7,
  407.9,
  404.9,
  369.8,
  366.5,
  363.6,
  360,
  350.5,
  414.6,
  409.3,
  406.4,
  405.7,
  394,
  402.7,
  402.2,
  397.9,
  375.5,
  382.3,
  379.3,
  373.3,
  349.6,
  343.1,
  338.3,
  336.7,
  338.6,
  360.5,
  370.4,
  385.1,
  385.4,
  385.3,
  364.2,
  353.5,
  327.4,
  329.4,
  345.5,
  357.8,
  382.6,
  376.4,
  372.2,
  367.1,
  378.8,
  375.7,
  383.2,
  373.4,
  369.3,
  383.4,
  390.6,
  379.7,
  364.2,
  361.4,
  376.4,
  385.6,
  382.3,
  357.7,
  346.6,
  341.8,
  388.8,
  350.3,
  337.1,
  337.1,
  335.3,
  333.7,
  335.9,
  337.9,
  338.7,
  337.4,
  338,
  341.1,
  342.1,
  346.5,
  344.6,
  340.7,
  355.9,
  355.4,
  350.3,
  353.7,
  359,
  357.5,
  362.4,
  365.7,
  375.5,
  325.1,
  314.8,
  358.6,
  355.3,
  361.7,
  381.1,
  394.7,
  377.5,
  366.5,
  376.9,
  378.1,
  375.6,
  377.8,
  380.2,
  385.2,
  385.2,
  382.8,
  376.5,
  368.8,
  393.8,
  391.7,
  377.7,
  362.6,
  395,
  368.9,
  358.5,
  355.2,
  354.2,
  352.3,
  355.2,
  358.4,
  356.4,
  356.3,
  363.6,
  368,
  351.6,
  352.3,
  361.3,
  349.4,
  347.5,
  353.3,
  345.8,
  343.8,
  342.8,
  342,
  339.2,
  338.6,
  338,
  339.2,
  343.1,
  349.4,
  359.2,
  365.5,
  370,
  375.1,
  391.9,
  397.4,
  380.4,
  382.4,
  395.5,
  390.5,
  388.9,
  392.8,
  394.9,
  407.4,
  406.1,
  409.6,
  399.5,
  403.4,
  391.3,
  389.4,
  411,
  379.6,
  374,
  373.3,
  369.8,
  363.6,
  366.1,
  369,
  370.7,
  367.2,
  365.5,
  364.9,
  356.9,
  359.4,
  361.3,
  361.4,
  360.1,
  359.4,
  359.7,
  360.2,
  357.1,
  357.3,
  355.2,
  351,
  345.3,
  347.3,
  353,
  357.5,
  364.6,
  367.2,
  366.9,
  370.6,
  369.8,
  371,
  367.5,
  363.6,
  371,
  372.8,
  374.9,
  370.7,
  369.7,
  368.5,
  370.9,
  368.3,
  361.3,
  361,
  363.5,
  363,
  403.6,
  379.4,
  378,
  377.4,
  372.9,
  369,
  364.2,
  359.1,
  351.2,
  347.2,
  344.6,
  341.5,
  339.9,
  338.9,
  339.5,
  337.7,
  337.6,
  336,
  333.2,
  329.6,
  331.8,
  324.9,
  313.6,
  312.4,
  316.1,
  324.1,
  329,
  331.4,
  336.9,
  342,
  342.6,
  348.9,
  350.1,
  352.7,
  352.3,
  349.2,
  354.6,
  358.4,
  359.3,
  361.9,
  368,
  365.6,
  365.8,
  358,
  355.9,
  357.6,
  349.6,
  346.4,
  407.9,
  401.8,
  393.2,
  375.8,
  344.6,
  344,
  346,
  346.5,
  348.9,
  352.1,
  347.8,
  352.1,
  349.3,
  345.8,
  344.3,
  364.1,
  378.9,
  377.2,
  379.5,
  371.6,
  356.7,
  342,
  335,
  332.2,
  329.6,
  331.4,
  336.3,
  343.6,
  352,
  360.5,
  362.2,
  362.1,
  366.9,
  371.7,
  386.6,
  381.5,
  385.5,
  384.9,
  395.2,
  388.6,
  383.2,
  399.4,
  378.3,
  380.8,
  384.6,
  373.8,
  370.6,
  372.4,
  403.1,
  384,
  380.5,
  378.3,
  373.1,
  371.8,
  370.7,
  370.5,
  364.5,
  366,
  366.5,
  369.1,
  362.2,
  363.3,
  366.7,
  365.7,
  362.9,
  359.3,
  358.3,
  356.3,
  354.4,
  356.3,
  356.5,
  356.1,
  353.7,
  355.6,
  356.8,
  357.9,
  361.5,
  365.6,
  370.6,
  373.8,
  376.3,
  380.7,
  392.6,
  389.5,
  386.2,
  382.6,
  384.3,
  381.7,
  379.9,
  377.8,
  376,
  373.9,
  371.9,
  371.4,
  373,
  438.6,
  391.6,
  383.7,
  390.4,
  396.2,
  397.2,
  400.5,
  388.6,
  386.9,
  391.7,
  390.1,
  386.8,
  381.2,
  382.3,
  397.8,
  401.4,
  406.8,
  411.6,
  414.2,
  406.9,
  410.6,
  405.2,
  402.3,
  397.1,
  396.7,
  394,
  397.5,
  403.1,
  404.6,
  413.5,
  419.4,
  419.9,
  420.6,
  420.1,
  423.8,
  423,
  423,
  421.2,
  419.6,
  419,
  417.8,
  417.1,
  417.9,
  418.3,
  419.2,
  419.8,
  419.7,
  420.1,
  429.4,
  423.1,
  420.4,
  418.9,
  418.4,
  417.7,
  417.7,
  417.3,
  417,
  417.3,
  417.3,
  417.3,
  417.1,
  416.7,
  416.1,
  415.7,
  415.8,
  415.3,
  415.1,
  415.1,
  415,
  415.1,
  414.9,
  415.3,
  415.2,
  415.5,
  415.8,
  417.6,
  418.9,
  422.7,
  424.4,
  433.4,
  439.7,
  445.3,
  447.7,
  429,
  428.6,
  427.6,
  426,
  427.8,
  422.9,
  421.4,
  419.9,
  419.7,
  419.8,
  422.6,
  422.6,
  421.1,
  455.4,
  427.9,
  401.5,
  384.9,
  383.5,
  380.5,
  377.6,
  376.5,
  377.5,
  377.9,
  377.6,
  376.8,
  376.7,
  375.5,
  375.6,
  375,
  381,
  389.4,
  379,
  383.4,
  381.6,
  371,
  371.1,
  371,
  366.7,
  364.5,
  369.4,
  379.8,
  395.5,
  400.1,
  404.1,
  397.6,
  392.5,
  394.2,
  397.1,
  393.8,
  390.9,
  398.5,
  400.7,
  400.8,
  400.1,
  397,
  399.3,
  399.5,
  405.7,
  394.6,
  390,
  389.3,
  445.3,
  406.4,
  392.7,
  394.3,
  388.3,
  383.3,
  383.7,
  384.4,
  387.1,
  399.6,
  398.6,
  406.7,
  419.7,
  416.4,
  416.5,
  417.5,
  416.9,
  417.8,
  416.4,
  415.6,
  414.2,
  413.3,
  414.1,
  414.5,
  417,
  420.1,
  424.4,
  425.9,
  432.1,
  410.8,
  393.4,
  389.5,
  393.5,
  396.9,
  397.9,
  396.6,
  395.4,
  403.1,
  429.6,
  407.8,
  416.3,
  416.4,
  419.3,
  434.6,
  416.3,
  409.8,
  412.8,
  408.3,
  416.5,
  409.9,
  392.9,
  403.1,
  409.8,
  396.5,
  400.9,
  389.4,
  388,
  390.1,
  396.5,
  401.8,
  405.8,
  407.8,
  404.1,
  400.5,
  397.8,
  398.2,
  403.2,
  406.2,
  406.4,
  405.4,
  407.1,
  403.6,
  404.4,
  407,
  408.7,
  415,
  422.2,
  428.8,
  431.7,
  397.6,
  399.8,
  388.6,
  406.8,
  405.5,
  407.2,
  397,
  400.4,
  399.3,
  397.2,
  398.6,
  399.1,
  403.6,
  394.9,
  392.3,
  383.7,
  372.8,
  440.3,
  365.8,
  345.4,
  343.5,
  342.3,
  350,
  361.9,
  371.3,
  379.7,
  386.2,
  385.9,
  382.9,
  375.6,
  377.4,
  381.7,
  378,
  385.2,
  388.1,
  390.8,
  388,
  387.5,
  391.1,
  392.9,
  394.7,
  396.5,
  398.8,
  402.1,
  403.1,
  404.3,
  401.7,
  390.9,
  373.3,
  366.4,
  377.2,
  392.3,
  374.7,
  372.9,
  385.7,
  391.8,
  391.9,
  395.1,
  393.9,
  407,
  407.2,
  399,
  396.1,
  397.6,
  403.2,
  417.4,
  407.8,
  403.3,
  402.1,
  391,
  390,
  392.9,
  389.9,
  380.7,
  369.6,
  374.7,
  377,
  381.1,
  388.8,
  393.9,
  397.6,
  399.6,
  399.1,
  395.5,
  397.3,
  402.5,
  401.5,
  400,
  397.4,
  400.9,
  400.7,
  402.2,
  403.6,
  405.8,
  406,
  406.3,
  407.4,
  405.4,
  403.9,
  407.6,
  410.5,
  414.3,
  401.8,
  392.5,
  389.9,
  382.1,
  362.4,
  358.6,
  377.8,
  356.8,
  351.9,
  349.2,
  359.6,
  386,
  360,
  340.2,
  341.1,
  336.8,
  319.2,
  315.3,
  316.7,
  329,
  345.4,
  317.1,
  312.8,
  312.8,
  330.6,
  333.6,
  378.6,
  376.1,
  363.4,
  358.9,
  350.1,
  371,
  364.8,
  352.5,
  352.2,
  333.7,
  337.5,
  344.6,
  362.2,
  371.3,
  379.1,
  373.6,
  376.8,
  381.9,
  384.2,
  375.9,
  382.9,
  379.5,
  374.1,
  361.6,
  362.8,
  365.7,
  368.1,
  341.4,
  331.1,
  353.8,
  340.5,
  338.1,
  338.6,
  374.4,
  362.8,
  336.2,
  320.6,
  314.5,
  313.6,
  310.5,
  308.6,
  308.5,
  308.3,
  308.9,
  308.5,
  306.3,
  304.9,
  300.8,
  306.2,
  317.9,
  322.6,
  323.9,
  325.7,
  336,
  345.5,
  344.7,
  348.6,
  350.3,
  356.6,
  359,
  371.2,
  373.2,
  371.2,
  372.3,
  377.6,
  382.3,
  386.7,
  388.2,
  387.7,
  388.9,
  393.6,
  395.6,
  395.9,
  396.4,
  396,
  395.3,
  394.8,
  394.4,
  394.4,
  398.7,
  402.2,
  447.7,
  409.8,
  400.8,
  400.3,
  401.5,
  400.7,
  399.8,
  402,
  403.1,
  402.6,
  395.7,
  395.7,
  392.8,
  340,
  357.3,
  387.1,
  388.1,
  386.6,
  384.3,
  383.5,
  384.7,
  383.4,
  383.7,
  380,
  384.4,
  379.1,
  378.6,
  373,
  340.9,
  345.7,
  361,
  347.1,
  357.3,
  367.9,
  361.1,
  369.4,
  363.7,
  372.2,
  366.4,
  365.7,
  358.1,
  367.5,
  385.4,
  372.8,
  370.4,
  358.1,
  361.4,
  360.4,
  385.9,
  365.3,
  365.4,
  352.9,
  352.6,
  352.2,
  352.6,
  351.8,
  353.9,
  358.8,
  361.4,
  359.3,
  358.9,
  359,
  361.8,
  364.5,
  359,
  360.5,
  360.9,
  371.9,
  359.1,
  349.4,
  344.9,
  342.9,
  337.5,
  333.7,
  335.7,
  336.6,
  343.1,
  351,
  356.8,
  366.8,
  356.2,
  354.2,
  356.4,
  352.5,
  348,
  357.3,
  355.7,
  352.9,
  355.3,
  347.7,
  349.3,
  378.9,
  379,
  384.9,
  362.6,
  375.1,
  390.1,
  384.1,
  377.8,
  388.1,
  397.7,
  396.1,
  395.8,
  394.9,
  392.2,
  389.4,
  388.4,
  389.7,
  388.6,
  386.7,
  385.8,
  384.7,
  381.6,
  380.4,
  378.7,
  378.2,
  378.6,
  379.2,
  379.8,
  380.7,
  381.6,
  384,
  386.1,
  391.5,
  394.3,
  401.5,
  404.9,
  405,
  411.9,
  420.5,
  373.8,
  365,
  338.4,
  361.3,
  368,
  367.6,
  361.5,
  346.5,
  357,
  356.4,
  346.3,
  344.5,
  346.6,
  370.3,
  394.1,
  348.1,
  327.5,
  321.8,
  321.8,
  321.7,
  323.8,
  324.1,
  323.6,
  322.1,
  322,
  322.3,
  318,
  317.4,
  316.4,
  316.8,
  312.4,
  315.4,
  316.9,
  321.6,
  324.9,
  336.7,
  336.8,
  338.7,
  322.5,
  297.1,
  289.4,
  301.5,
  310.9,
  315,
  320.8,
  329.5,
  340.5,
  355.1,
  349.7,
  347.7,
  338.2,
  345.3,
  356.9,
  360,
  351.2,
  341.6,
  339.7,
  342.9,
  336,
  336,
  338.6,
  340.4,
  370.9,
  353.5,
  356.2,
  358.4,
  362.5,
  364.1,
  375,
  374.9,
  374.1,
  375.8,
  375.4,
  383.6,
  388.2,
  385.6,
  380.3,
  378,
  378.9,
  377,
  381.7,
  390,
  392.2,
  390.4,
  390.5,
  390.4,
  389.2,
  391.9,
  387.9,
  372.3,
  379.1,
  382,
  383.5,
  374.2,
  380.2,
  389.7,
  385.5,
  380.6,
  392.1,
  389.1,
  383.7,
  360.6,
  367.5,
  398.7,
  400.6,
  383.4,
  386.5,
  403.5,
  397.2,
  431.3,
  399.4,
  365.5,
  350,
  349.4,
  348.9,
  344.9,
  366.5,
  387.9,
  394,
  388.8,
  379.5,
  360.7,
  364.6,
  381.9,
  382.6,
  359.7,
  335,
  336.4,
  340.1,
  365.1,
  347.4,
  381.3,
  371.2,
  375.2,
  381.9,
  381.3,
  382.8,
  377.1,
  361,
  346.3,
  347.4,
  373.9,
  385.4,
  374,
  374.4,
  369.7,
  368.2,
  361.3,
  349.5,
  355,
  346.7,
  350,
  357.2,
  383.2,
  373.6,
  373.6,
  369.6,
  388.4,
  383.2,
  380.1,
  369.1,
  361.9,
  353.2,
  327.5,
  316.1,
  316.1,
  312.7,
  311.7,
  309.3,
  310.4,
  315.9,
  312.5,
  320.8,
  313.4,
  308.2,
  310.7,
  342.2,
  361.5,
  354.5,
  365,
  342.5,
  310.9,
  308.1,
  304.9,
  348.6,
  316.8,
  308.9,
  321.4,
  353.9,
  351.8,
  357.2,
  326.9,
  344.9,
  340.2,
  335,
  344.9,
  346.8,
  335.3,
  329.9,
  330.4,
  339.5,
  320.9,
  313.1,
  310.3,
  308.7,
  396.5,
  327.9,
  309.8,
  344.9,
  320.4,
  309.4,
  310.2,
  313.5,
  324,
  331,
  354.2,
  371.7,
  374.7,
  383.4,
  382.1,
  382,
  382.5,
  382.2,
  382.6,
  382.2,
  382.4,
  382.7,
  383.4,
  383,
  383.4,
  382.7,
  384.1,
  385.4,
  388,
  389.4,
  391.9,
  396.6,
  396.4,
  402.4,
  402,
  390.8,
  374.2,
  377.9,
  376.3,
  367.7,
  369.3,
  371.5,
  379.5,
  341.5,
  332.3,
  333,
  362.4,
  345.8,
  392,
  350,
  322.2,
  324,
  339.1,
  330.3,
  325,
  320.9,
  318,
  323.4,
  337.6,
  346.8,
  351.5,
  363.3,
  358.7,
  360.6,
  363.1,
  367.4,
  368.6,
  376.9,
  375.9,
  374,
  372.3,
  378.3,
  374.6,
  383.5,
  384.1,
  386.7,
  383.7,
  342.2,
  350.8,
  352.8,
  361.6,
  376,
  382.3,
  381.2,
  376.4,
  364.5,
  369,
  367.1,
  371.9,
  346.9,
  378.3,
  379.1,
  382.4,
  385.2,
  386.8,
  385.9,
  389,
  385.9,
  376,
  367.4,
  370.6,
  374.5,
  376,
  370.4,
  368.6,
  375,
  337.9,
  343.9,
  356.9,
  379.6,
  364.5,
  329.9,
  338.8,
  347.2,
  343.2,
  316,
  307.2,
  328.5,
  337.4,
  362,
  358.3,
  369.6,
  368.7,
  367.6,
  368.1,
  362.6,
  360,
  370.4,
  360.4,
  365.6,
  348.7,
  361.6,
  340.9,
  350.5,
  349.2,
  347,
  334.2,
  351.6,
  363.9,
  353.6,
  328.4,
  325,
  303.9,
  301.4,
  381.7,
  312.4,
  344,
  342.3,
  289.2,
  290.7,
  297.6,
  309.4,
  348.7,
  344.7,
  334,
  356.7,
  356.8,
  355.9,
  353.3,
  350.9,
  353.3,
  353.6,
  349.5,
  334.3,
  332.3,
  320.8,
  338.7,
  354.3,
  349.4,
  335.6,
  345.7,
  317.1,
  339.2,
  327.8,
  298.4,
  336.6,
  351.1,
  344,
  359.3,
  361.3,
  363.2,
  348.5,
  348.3,
  341.5,
  349.2,
  333.4,
  353,
  355.6,
  345.9,
  319.1,
  309.6,
  308.4,
  375.1,
  323.1,
  309.9,
  310.4,
  311,
  310,
  311.5,
  312.4,
  312.2,
  314.7,
  314.3,
  311.2,
  304.6,
  304.8,
  305,
  304.1,
  302.7,
  303.1,
  304.4,
  306.9,
  307.2,
  308.2,
  323.6,
  312.2,
  317.1,
  315.6,
  308.5,
  304.5,
  301.3,
  304.4,
  308,
  322.4,
  335.4,
  330.8,
  342.6,
  347.3,
  354.3,
  357.8,
  356.3,
  361.8,
  358.2,
  359,
  353.3,
  352.8,
  353.2,
  367.3,
  369.5,
  355.1,
  397.4,
  331.1,
  315.2,
  317.4,
  321.7,
  316.3,
  317.9,
  321.8,
  325.1,
  325.9,
  326.6,
  330.8,
  331.6,
  344.7,
  333.6,
  343.2,
  359.6,
  366.4,
  364.5,
  380,
  385,
  385.2,
  385.9,
  387.1,
  387.7,
  375.9,
  366.6,
  370,
  370.1,
  370,
  367.6,
  361.5,
  356.5,
  339.9,
  330.4,
  340.5,
  337.7,
  374.3,
  365.1,
  346.8,
  366.9,
  380.1,
  383.1,
  385,
  374.7,
  376.1,
  379.9,
  379.4,
  411.8,
  375.3,
  347.1,
  377.9,
  377.4,
  370.1,
  379.9,
  379.4,
  377.7,
  378.5,
  378.1,
  377.1,
  374.9,
  373.4,
  372.6,
  373.5,
  364.1,
  368.3,
  369.8,
  366.5,
  364,
  358.3,
  352.6,
  349.2,
  348.5,
  345.7,
  323.3,
  288.3,
  319.3,
  288.2,
  294,
  313.3,
  315.6,
  303.5,
  310.1,
  303,
  298.2,
  299.8,
  299.1,
  303.2,
  299.9,
  333.5,
  321.3,
  330.1,
  340.9,
  290.9,
  328.2,
  295.2,
  330.4,
  330,
  310.1,
  298.6,
  335,
  322.4,
  296.2,
  294.3,
  334.7,
  349.2,
  329.5,
  311.4,
  309.4,
  308.6,
  307.8,
  318.5,
  344.9,
  331.7,
  324.7,
  344.4,
  344.3,
  341.5,
  329.2,
  324.9,
  333.3,
  343.4,
  328.5,
  329.1,
  310.9,
  285.8,
  290.2,
  297.7,
  321.3,
  312.5,
  331,
  328,
  323.2,
  321.4,
  317.8,
  336.7,
  348.7,
  334.7,
  312.9,
  310.6,
  315.3,
  316.5,
  335.3,
  342.3,
  332.9,
  312.6,
  299.3,
  297.1,
  296.3,
  297.8,
  310.4,
  294.7,
  295.8,
  295.6,
  295,
  293.1,
  292.4,
  292.6,
  311,
  294.8,
  292.2,
  292.6,
  290.6,
  294.5,
  302.2,
  309.6,
  323.1,
  327.3,
  294.4,
  290.9,
  286.2,
  285.1,
  285.6,
  288.8,
  296.9,
  308,
  315.9,
  313.9,
  315.3,
  317.3,
  320.6,
  316,
  326.1,
  334.6,
  331,
  325.8,
  333.6,
  318.8,
  319,
  326.3,
  332.3,
  320.6,
  349.1,
  314.9,
  309.3,
  314.1,
  306.7,
  305.8,
  301.9,
  303.3,
  311.2,
  311.5,
  300.1,
  314.2,
  327.2,
  328.1,
  310.9,
  304.3,
  311.2,
  314.3,
  336.5,
  329.2,
  304.2,
  306.8,
  292.4,
  290,
  285.4,
  281.6,
  280.7,
  285.2,
  287,
  291.9,
  298.6,
  303.5,
  305.6,
  308,
  314.5,
  312.7,
  314,
  312.2,
  317.1,
  318.9,
  319.9,
  319.7,
  319.6,
  317.1,
  317.2,
  320.6,
  322.4,
  385,
  355.8,
  336,
  338.4,
  344.4,
  336.3,
  325.4,
  322.5,
  321.5,
  319.3,
  317.5,
  323.6,
  317.5,
  310.4,
  308.1,
  307.1,
  306.2,
  304.8,
  304.9,
  304,
  306.5,
  304.1,
  311.4,
  313.1,
  310.8,
  309.2,
  303.8,
  297.8,
  297.5,
  303.3,
  309.3,
  320,
  321.6,
  334.1,
  358.1,
  384.8,
  392,
  393.3,
  393.9,
  392.6,
  393.4,
  392.1,
  393.8,
  394.5,
  392.8,
  393.2,
  390.1,
  388.9,
  421.3,
  402.5,
  389.4,
  387.2,
  386.2,
  385.8,
  384.4,
  365.2,
  351.6,
  332.2,
  327.4,
  325.3,
  325.2,
  325.7,
  325.6,
  327,
  335.4,
  336.4,
  321.8,
  320.9,
  320.1,
  323.8,
  345.7,
  351.9,
  352.4,
  359.3,
  367.9,
  367.4,
  356.8,
  350.9,
  325.7,
  357.5,
  373.5,
  373.6,
  352.3,
  383,
  373.6,
  337.5,
  335.9,
  342.3,
  346.5,
  358.6,
  356.1,
  367.7,
  349.8,
  344.2,
  337.9,
  366.7,
  404.5,
  349.9,
  330.9,
  323.8,
  315.4,
  319.7,
  313.5,
  314.4,
  315.5,
  310.8,
  312.2,
  331.4,
  333.5,
  346.9,
  348.5,
  353.7,
  357.1,
  358.6,
  359.1,
  356.7,
  356.5,
  355.6,
  337.7,
  334.2,
  345.1,
  334,
  328.7,
  350.8,
  345.3,
  326.6,
  316.1,
  314.8,
  310,
  310.5,
  317,
  316.1,
  317.3,
  328.5,
  335.1,
  333.1,
  355,
  340.1,
  320.1,
  328.3,
  317,
  320.4,
  297.6,
  287.9,
  357.9,
  308.2,
  292.4,
  289.2,
  284.1,
  280.7,
  280.8,
  282.7,
  284.1,
  282.5,
  279.2,
  279,
  277,
  278.7,
  277.4,
  278.2,
  277.1,
  275.9,
  276.5,
  276.2,
  279,
  280.1,
  279.3,
  277.4,
  277.6,
  285.2,
  259.9,
  246.1,
  255.9,
  270.5,
  274.4,
  279.1,
  284.2,
  288.3,
  302.4,
  297.2,
  301.2,
  302,
  305.9,
  305.5,
  309.4,
  304.1,
  307.8,
  291.6,
  299.5,
  288.3,
  287.3,
  294,
  325.7,
  303.4,
  288.6,
  288.2,
  285.7,
  286.1,
  283.7,
  284.1,
  286.3,
  283,
  282.4,
  280.9,
  278.2,
  277.6,
  277.1,
  276.1,
  275.4,
  276.1,
  275.8,
  275.2,
  274.7,
  273.8,
  273.7,
  273.9,
  273.8,
  273.3,
  270.2,
  268.7,
  270.9,
  275.6,
  277.7,
  281.1,
  284.1,
  289.3,
  293,
  296.2,
  295.9,
  296.1,
  296.6,
  299.8,
  300.7,
  300,
  299.5,
  298.3,
  295.8,
  295.7,
  293.3,
  291.7,
  370.4,
  314,
  297.7,
  296.2,
  293.7,
  293.9,
  292.9,
  290.7,
  288.5,
  286.1,
  283.9,
  283.1,
  282.5,
  281.3,
  281.3,
  280.2,
  279,
  278.5,
  277.9,
  277.1,
  277.3,
  275.3,
  274.5,
  274.6,
  274.3,
  273.8,
  270.3,
  268.4,
  270,
  272.5,
  276.5,
  281.2,
  286.7,
  292,
  296.4,
  298.7,
  300.9,
  297.3,
  300,
  306.7,
  308,
  310.6,
  310.6,
  308.1,
  306.9,
  304.6,
  302.5,
  300.3,
  372,
  317.7,
  302.3,
  301.6,
  299.1,
  297.1,
  296,
  294.5,
  290.5,
  288,
  287.7,
  285.7,
  285.5,
  285.7,
  286.4,
  286.4,
  286.6,
  285.4,
  284.7,
  284.6,
  283.6,
  283.4,
  285.3,
  285.2,
  286.2,
  285.9,
  282.2,
  279.2,
  278.1,
  280.8,
  286.2,
  288.5,
  307.8,
  323.5,
  331.9,
  318.8,
  313.7,
  309.8,
  310,
  310.3,
  313.4,
  318.5,
  323.8,
  337.1,
  361.4,
  374.1,
  366.5,
  346.1,
  386.5,
  373.9,
  364.6,
  341.5,
  360.1,
  369.8,
  369.8,
  369.3,
  369.9,
  349.2,
  319.2,
  314.8,
  312.1,
  309.9,
  314.1,
  309.3,
  311.7,
  355,
  362.8,
  364.4,
  364.2,
  365.1,
  365.6,
  366.2,
  367.6,
  367.7,
  368.5,
  368.4,
  368.3,
  368.1,
  368.7,
  370.3,
  371.6,
  373.2,
  374.7,
  378.7,
  379.7,
  380.8,
  379.1,
  380.5,
  381.2,
  380.5,
  380.9,
  380.1,
  379.5,
  378.6,
  379.1,
  378.4,
  394.7,
  379.4,
  372.1,
  365.5,
  366.3,
  369.3,
  344.4,
  307.4,
  305.4,
  302.9,
  301.1,
  299.6,
  301.4,
  300.5,
  298.6,
  297.1,
  297.3,
  297.1,
  297.6,
  299.3,
  300,
  298.4,
  297.5,
  298.1,
  296.1,
  295,
  290.9,
  286.6,
  287.7,
  291.5,
  294.6,
  298.3,
  306.1,
  311.6,
  316.1,
  321,
  321.8,
  316.6,
  319,
  325,
  324.8,
  325.8,
  326.3,
  325.8,
  324.7,
  324,
  321.7,
  321,
  377.2,
  331.6,
  319.8,
  319.5,
  312.5,
  317.9,
  313.1,
  310.4,
  307,
  308.3,
  307.7,
  309.1,
  306,
  304.7,
  304.8,
  303.3,
  301.8,
  302.1,
  299.9,
  300.6,
  302.6,
  301.6,
  296.5,
  295.6,
  297.4,
  294.7,
  291.8,
  287.4,
  288.6,
  292.4,
  294.3,
  298.1,
  301.8,
  306,
  311.9,
  315.8,
  319.4,
  317.9,
  322,
  329.6,
  331.6,
  331.9,
  331.2,
  330.2,
  328.7,
  326.8,
  323.3,
  319.2,
  372.2,
  329.2,
  321.3,
  315,
  307.2,
  304.9,
  302.2,
  300.3,
  298.9,
  297.6,
  296.3,
  294.4,
  293,
  292.3,
  292.1,
  321.1,
  366.4,
  367.7,
  366.7,
  365.8,
  365.5,
  365.9,
  366.2,
  366.6,
  365.9,
  366.5,
  366.1,
  366.2,
  366.7,
  367.2,
  367.7,
  367.2,
  367.6,
  368,
  368.1,
  368.2,
  368.1,
  368.3,
  364.3,
  339.6,
  322.3,
  305.3,
  304.5,
  305.6,
  304.2,
  302.2,
  303.6,
  304.1,
  354.5,
  319.1,
  311.1,
  300.2,
  295.8,
  291,
  288.7,
  289.8,
  290.2,
  288.6,
  289.2,
  289.4,
  286.4,
  287.2,
  292.1,
  294.5,
  287.5,
  292.5,
  302.7,
  309.4,
  326.5,
  336.8,
  339,
  339.8,
  340.1,
  340.6,
  340.7,
  339.3,
  339,
  340.6,
  345.9,
  342,
  347.4,
  352,
  351.8,
  317.2,
  290.8,
  293.7,
  310.2,
  315.7,
  310.9,
  312.9,
  313,
  311.6,
  310.9,
  309,
  305.7,
  303.9,
  335.4,
  304.4,
  307,
  310,
  311.3,
  316.9,
  314.5,
  315.4,
  310.4,
  301.7,
  315.7,
  311.9,
  304.9,
  331.4,
  331,
  329.2,
  322.9,
  324.1,
  323.3,
  332.9,
  333.9,
  333.1,
  332.6,
  330.9,
  330.6,
  335,
  336.3,
  333.4,
  333.9,
  342.7,
  349.9,
  356,
  361.8,
  357.7,
  336.6,
  332.3,
  339.8,
  344.2,
  343.8,
  361.1,
  360.4,
  333.8,
  343.2,
  356,
  349.9,
  348.9,
  355,
  412,
  373.4,
  359.1,
  375.7,
  369.1,
  363.8,
  372.4,
  370.2,
  366.8,
  366,
  367.7,
  377.9,
  374.6,
  376,
  377.5,
  380.9,
  379.1,
  378.4,
  379,
  377.8,
  381,
  382.8,
  384,
  383.8,
  385,
  386.1,
  386.4,
  386.1,
  384.6,
  386.3,
  387.8,
  388.1,
  389.4,
  387.5,
  381.7,
  373.9,
  377,
  375,
  378.3,
  375,
  373.8,
  370.2,
  384.8,
  380.6,
  386.9,
  382.4,
  386,
  387.4,
  406.4,
  392.7,
  388.4,
  392.4,
  393.3,
  392.3,
  396.2,
  396.8,
  392.8,
  389.6,
  387.6,
  386.1,
  385,
  384.4,
  384.7,
  385.2,
  385.3,
  385.3,
  386.1,
  386.2,
  386.2,
  386.3,
  387.1,
  387.2,
  387.7,
  388.3,
  388.5,
  389.3,
  391.1,
  394.1,
  397.6,
  400.7,
  402.4,
  403.2,
  405.8,
  406.7,
  406.1,
  403.3,
  402,
  402.2,
  403.9,
  403.8,
  404.1,
  401.4,
  399.6,
  400.4,
  399.9,
  397.5,
  410.4,
  400.9,
  396.2,
  372.1,
  376.2,
  377.6,
  386.6,
  389.1,
  391.2,
  363.3,
  373.7,
  382.7,
  377.2,
  376.2,
  376.7,
  372.8,
  372.8,
  369.2,
  358.1,
  346.8,
  347.1,
  352.8,
  368.6,
  367.4,
  367.1,
  366.7,
  367,
  365.4,
  364.1,
  353.6,
  334.3,
  342.1,
  331.6,
  335.7,
  362.5,
  348.2,
  359.8,
  363.7,
  300.4,
  313.8,
  353,
  307.8,
  331.2,
  359,
  358.1,
  354.7,
  363,
  353.3,
  396.1,
  362.8,
  347.9,
  354.9,
  321.5,
  329.6,
  306.6,
  285.3,
  282.7,
  337.6,
  321.9,
  344,
  349.5,
  343.6,
  346.2,
  317.5,
  283.3,
  286.7,
  289.8,
  300.9,
  299.3,
  296,
  290.7,
  296,
  315.9,
  297.8,
  300.3,
  316.6,
  319.2,
  326.3,
  295.3,
  292.6,
  307.7,
  333.6,
  333.4,
  345.2,
  361.5,
  361.6,
  368.9,
  362.5,
  363.2,
  360.6,
  368.9,
  366.5,
  364.2,
  361.4,
  363.8,
  362.9,
  393.9,
  348.6,
  362.6,
  341,
  338.9,
  346.6,
  367.3,
  317.8,
  298.3,
  312.4,
  350.1,
  363,
  362.5,
  364.7,
  368.6,
  366.3,
  365.4,
  368.2,
  366.2,
  365.7,
  369.2,
  371.5,
  369.2,
  367.8,
  366.7,
  369.4,
  368.9,
  364.2,
  364.8,
  368.7,
  369.7,
  367.5,
  356.8,
  354.7,
  366.7,
  345.9,
  376.8,
  382,
  382.5,
  383.4,
  383.3,
  382.7,
  382.3,
  381.7,
  382.4,
  382.1,
  382.8,
  382.5,
  399,
  386.4,
  379.6,
  378.4,
  365.1,
  317.1,
  312.8,
  312.4,
  310.6,
  310.9,
  311.4,
  311.1,
  312.2,
  312.2,
  311.9,
  311.5,
  311.4,
  312,
  312.2,
  313.7,
  346.9,
  363.4,
  375.1,
  375.3,
  377.6,
  378.3,
  378.6,
  379.9,
  379.4,
  378.7,
  378.3,
  377.2,
  376,
  376.9,
  377,
  377.3,
  377.4,
  377.9,
  378.7,
  379.4,
  379.6,
  380,
  384.1,
  384.3,
  382.2,
  382.9,
  379,
  379.8,
  384.1,
  378,
  374.4,
  374.6,
  373.9,
  373.1,
  370.8,
  370.5,
  372.7,
  372.5,
  372.6,
  373.1,
  372.5,
  371.8,
  371.7,
  371,
  369.6,
  367.8,
  363,
  356.8,
  335.4,
  306.8,
  297.3,
  295.5,
  294.8,
  313.2,
  313.1,
  295.3,
  294.9,
  294,
  296,
  300.6,
  305.4,
  303,
  303,
  304.8,
  308.6,
  312.1,
  308.1,
  313.2,
  317.9,
  322.7,
  332.1,
  343.5,
  336.8,
  331.4,
  334.6,
  339.9,
  378.7,
  362,
  353.5,
  346.9,
  343.8,
  349.3,
  347.3,
  345.2,
  351.5,
  350.8,
  351.7,
  345.8,
  348.1,
  362.2,
  373.3,
  390.4,
  395,
  400.8,
  398.7,
  399.7,
  398.8,
  398,
  397.6,
  397.4,
  398.2,
  397.9,
  397.9,
  398.9,
  399.5,
  399,
  399.5,
  400.2,
  400.4,
  401,
  398,
  397.6,
  383.2,
  380.8,
  355.1,
  389,
  378.7,
  386.2,
  369,
  344.1,
  376.9,
  375.2,
  374.1,
  373.7,
  404.5,
  327.5,
  299.7,
  312,
  319.1,
  310,
  297.9,
  309.5,
  297.7,
  296.2,
  302.4,
  300.3,
  295.9,
  317.9,
  311.6,
  315.3,
  308.2,
  304.6,
  318.7,
  315.6,
  340,
  344.7,
  335.5,
  351.1,
  350.5,
  347.3,
  330.8,
  331.5,
  318.3,
  323.6,
  346.8,
  371.1,
  377.2,
  378,
  380.6,
  383.7,
  385,
  386.9,
  388.8,
  391,
  393.1,
  390.1,
  393.2,
  393.2,
  394.3,
  396.5,
  397.1,
  397.1,
  408.4,
  389,
  391.4,
  390.7,
  390.2,
  391.2,
  392.6,
  393.5,
  394.6,
  396.6,
  398.1,
  399.2,
  400,
  401.2,
  401.7,
  398.9,
  393.3,
  387.5,
  400.7,
  402.9,
  403.3,
  402.6,
  401,
  400.7,
  401.1,
  399.3,
  399.9,
  399.9,
  400.9,
  401.4,
  393.9,
  394.8,
  372.5,
  363.1,
  392.8,
  391.9,
  390.1,
  390.8,
  390.5,
  393.3,
  394.8,
  392.2,
  389.8,
  391.1,
  387.8,
  389.3,
  387.1,
  384.2,
  380.8,
  377.1,
  383.4,
  383.5,
  388.3,
  375.8,
  384.2,
  384.6,
  384,
  384.2,
  380.9,
  384.7,
  386.2,
  385.5,
  384.4,
  393.4,
  393.2,
  390.1,
  390.1,
  389.6,
  389.1,
  391.3,
  389.8,
  390,
  383.1,
  373.6,
  385.8,
  388.6,
  379.9,
  365.7,
  318.1,
  306.8,
  305.7,
  295.9,
  320,
  341.7,
  337.3,
  353.9,
  353.5,
  362.4,
  348.9,
  349.5,
  344,
  332,
  325.8,
  307.5,
  331.6,
  314.8,
  353.4,
  340,
  369.2,
  368.9,
  363,
  367.3,
  318.9,
  333.9,
  352.3,
  365.5,
  367.2,
  367.9,
  363.9,
  359.5,
  363.1,
  362.6,
  366.3,
  359.7,
  367.3,
  359.5,
  342.2,
  351.5,
  333.6,
  303.6,
  332.4,
  289.4,
  288.3,
  322.5,
  317,
  339.3,
  363.6,
  368,
  369.6,
  372.2,
  369.5,
  343.5,
  338,
  326.5,
  325.7,
  315.7,
  316.2,
  322.8,
  340,
  350.9,
  346.6,
  327,
  333.1,
  339.1,
  351,
  343.1,
  352.3,
  341.4,
  342.3,
  345.1,
  342.6,
  355.6,
  365,
  363.9,
  362.6,
  361.7,
  360.8,
  360.8,
  361,
  360.4,
  360.3,
  359.6,
  359.1,
  356.8,
  354.5,
  350.7,
  348,
  347.1,
  344.1,
  341.5,
  343,
  342.3,
  342.5,
  341.4,
  344.9,
  364.8,
  372,
  382.3,
  347.3,
  340.5,
  350.4,
  361.4,
  366,
  343.2,
  282.2,
  291.7,
  326.4,
  353.5,
  310,
  313.8,
  304.4,
  354,
  316.7,
  324.2,
  350,
  337.2,
  347.9,
  348.1,
  345.6,
  348.4,
  342.5,
  334.5,
  334.6,
  331.2,
  328,
  328.1,
  327.3,
  326.2,
  327.8,
  329.7,
  337,
  346.3,
  344.8,
  341.8,
  324.6,
  331.2,
  338.9,
  337.4,
  322.4,
  319.5,
  330.1,
  342.5,
  332.2,
  337.9,
  333.2,
  327.1,
  337.1,
  345.8,
  338,
  334,
  347.5,
  334.9,
  329.1,
  332.7,
  340.3,
  328,
  311.8,
  292.3,
  308.1,
  415.3,
  340.4,
  348.7,
  336.3,
  339.2,
  348.1,
  349.1,
  322.7,
  330.3,
  341.5,
  344.2,
  333.8,
  350,
  351.8,
  352.2,
  349.7,
  343.8,
  310.4,
  319.8,
  312.3,
  332.6,
  321.4,
  303.7,
  318.2,
  310.6,
  284.3,
  296.4,
  302.1,
  331,
  326.2,
  309.7,
  295.9,
  348.7,
  340.7,
  347.6,
  283.5,
  347.2,
  344.5,
  308.1,
  291.8,
  309.3,
  311.9,
  345.3,
  348.8,
  332.1,
  333,
  336.6,
  338.3,
  364.8,
  347.7,
  332.9,
  337.6,
  345.6,
  346.9,
  350.1,
  352.2,
  352.6,
  352.6,
  352.9,
  352.6,
  352.1,
  352,
  352.7,
  352.6,
  352.4,
  352,
  352,
  352.1,
  351.4,
  351.4,
  351.5,
  351.5,
  351.6,
  351.8,
  350.9,
  350.5,
  349.6,
  349.3,
  349,
  346.4,
  344.4,
  344.3,
  346.3,
  346.9,
  346,
  348.4,
  348.2,
  347.9,
  347.9,
  347.8,
  340.2,
  312.7,
  316.8,
  323.5,
  345.3,
  345.5,
  346.5,
  313.6,
  284.9,
  287.6,
  303.5,
  285,
  297.5,
  306.3,
  324.2,
  345.1,
  335.9,
  337.9,
  340.6,
  346.1,
  344,
  341.5,
  340.5,
  329.4,
  333.7,
  339.2,
  341.5,
  340.4,
  336.3,
  335.1,
  336.4,
  337.8,
  337.5,
  338.7,
  339.3,
  340.3,
  341.2,
  342.3,
  342.1,
  342.4,
  342.9,
  342.6,
  342.2,
  339.2,
  318.1,
  294.4,
  324.2,
  335.2,
  338.3,
  325.8,
  329.3,
  329.9,
  335,
  325.4,
  353.9,
  341.9,
  310.1,
  321.7,
  326,
  335.4,
  341.1,
  341.3,
  342,
  344.8,
  346,
  343.3,
  342.6,
  347.8,
  346.4,
  347.8,
  352.2,
  354.1,
  355.5,
  357.3,
  358.8,
  359.5,
  360.5,
  362.6,
  363.4,
  363.7,
  363.5,
  363,
  363.5,
  363.5,
  364.2,
  365.4,
  367,
  369.4,
  370.6,
  369.8,
  370.4,
  370.1,
  371.4,
  373.2,
  363.9,
  375,
  371.7,
  380.5,
  379.5,
  380,
  380.4,
  371.4,
  397.7,
  335.1,
  316.4,
  318.1,
  316.4,
  312.8,
  309.5,
  308.3,
  309.2,
  305.1,
  303.1,
  301.2,
  299.8,
  298.6,
  296.7,
  296,
  295.8,
  295.8,
  295.7,
  294.9,
  294.1,
  293.2,
  292.5,
  292.8,
  291.8,
  292.1,
  291.3,
  290.3,
  290,
  288.8,
  286.7,
  285.8,
  287.2,
  291.2,
  296.8,
  300.8,
  304.6,
  307.1,
  309.3,
  305.7,
  311.7,
  317.3,
  319.1,
  320.1,
  320.5,
  320.8,
  321.6,
  321.1,
  391.4,
  344.4,
  323.7,
  320.4,
  318.6,
  317.8,
  317.1,
  318,
  315.5,
  311.8,
  312,
  311.9,
  311.1,
  311.5,
  311.5,
  310.6,
  308.6,
  308.2,
  306.9,
  308,
  313.2,
  308.2,
  308.1,
  311.5,
  313.4,
  313,
  308.4,
  304.9,
  304.5,
  301.6,
  295.4,
  294.6,
  291.1,
  292.5,
  298.4,
  304.2,
  305.6,
  307.5,
  309.8,
  309.2,
  314.6,
  320.7,
  326.3,
  327.6,
  327.3,
  327.5,
  328.8,
  326.3,
  379.9,
  341.9,
  332,
  329.3,
  330.7,
  330.3,
  328.7,
  327.3,
  326.1,
  320.7,
  319.4,
  319.3,
  322,
  316.3,
  327.2,
  371.5,
  370,
  370.4,
  376.8,
  377.4,
  377.9,
  377.4,
  376.8,
  373.4,
  367.2,
  371.6,
  372.3,
  368.7,
  362.8,
  365.9,
  366,
  362.4,
  357.7,
  356.2,
  355,
  354.5,
  353.7,
  354,
  353.4,
  351.7,
  350.3,
  344.1,
  306.8,
  286.5,
  276.5,
  282.6,
  283.3,
  270.4,
  301.6,
  268.1,
  258.9,
  260.9,
  257.1,
  258.2,
  263.2,
  267.7,
  278.3,
  288.1,
  276.4,
  277.4,
  287.6,
  286.3,
  281.2,
  263,
  251.7,
  245,
  242.5,
  240.5,
  244.3,
  245.7,
  246.3,
  247.6,
  247.9,
  247.2,
  244.3,
  251.5,
  269.2,
  274.9,
  267.7,
  244.2,
  231.8,
  235.3,
  243.8,
  271.4,
  294.8,
  262.6,
  248.4,
  243.1,
  249.7,
  254.9,
  256.4,
  254.9,
  255.2,
  254.7,
  256.9,
  257.4,
  311.8,
  274.2,
  263.7,
  257.4,
  255.5,
  251.8,
  247.8,
  244.6,
  247.6,
  244.9,
  243.2,
  242.1,
  241.9,
  241.5,
  241.6,
  242.9,
  244.8,
  240.7,
  240.9,
  242.2,
  239.7,
  239.3,
  240.3,
  239,
  238.6,
  237.8,
  239.2,
  236.6,
  237.2,
  238.1,
  229.6,
  225.8,
  228.6,
  231.4,
  233.2,
  237.3,
  242.4,
  242.2,
  245.6,
  239.1,
  245.3,
  248.9,
  251,
  250.8,
  253,
  251.9,
  252.9,
  250.6,
  316.7,
  272,
  259.1,
  267.3,
  270.6,
  268.8,
  264,
  267.3,
  269.1,
  271.1,
  270.2,
  275.2,
  333.8,
  342.1,
  338.1,
  335.4,
  304,
  283.8,
  269.6,
  270.3,
  281.9,
  329.6,
  336.6,
  341.3,
  340.3,
  332.3,
  341.6,
  335.7,
  335.3,
  337.6,
  335.6,
  334.4,
  332.6,
  331.2,
  331.1,
  331.7,
  334.4,
  334.8,
  320.9,
  315.3,
  346.8,
  339.7,
  338.5,
  307.5,
  333.8,
  340,
  288.5,
  332.1,
  346.6,
  322.5,
  280.2,
  333.5,
  304.4,
  316.2,
  323.6,
  327.8,
  304,
  312.6,
  280.7,
  322.5,
  317.7,
  306.5,
  344.2,
  343.8,
  343.3,
  342.7,
  342.6,
  334.1,
  332.9,
  331.2,
  323.9,
  327.7,
  328.1,
  323.3,
  306.4,
  297.3,
  311,
  305.8,
  279.1,
  257.1,
  289.8,
  296.8,
  316.9,
  316.6,
  285.6,
  292.4,
  297.5,
  306.5,
  286.6,
  311.4,
  288.3,
  299.6,
  294.4,
  283.5,
  262.7,
  282.3,
  336.6,
  330.5,
  312,
  305.5,
  285.9,
  282.2,
  294.3,
  297.3,
  296.7,
  287.2,
  304.1,
  313.4,
  326.8,
  322.6,
  312,
  274,
  277.7,
  264.8,
  262.6,
  291.8,
  269.8,
  279.2,
  290.5,
  295.4,
  295,
  306.6,
  301.4,
  321.4,
  321.9,
  328.8,
  331.9,
  334.7,
  335.3,
  337.3,
  340.1,
  341.6,
  337.1,
  344.7,
  346.7,
  339.4,
  337.1,
  327.7,
  347.7,
  348.5,
  350.1,
  344.9,
  348.4,
  350.9,
  355.4,
  353.3,
  353.2,
  352.9,
  352.1,
  351.9,
  351.9,
  350.9,
  348.5,
  347.7,
  346.9,
  347.5,
  345.2,
  344.9,
  343.7,
  324.1,
  316.8,
  308.7,
  306.6,
  315.5,
  339.8,
  334.3,
  318.9,
  317.9,
  323.3,
  332.9,
  336.9,
  337.6,
  337,
  336.8,
  335.1,
  330.2,
  327,
  322.4,
  290.2,
  277.1,
  294,
  313.1,
  307.9,
  328.2,
  334.2,
  345.1,
  347.5,
  349.9,
  345.3,
  348.4,
  345.2,
  371.1,
  352.5,
  343.5,
  345.4,
  345,
  350.2,
  349.1,
  350.6,
  348,
  345.6,
  342.2,
  339.7,
  338.9,
  333.1,
  329.9,
  324.4,
  319.2,
  319.3,
  326.2,
  324.1,
  327.8,
  325.6,
  322.8,
  317,
  298.4,
  269.3,
  252.2,
  244.5,
  241.9,
  240,
  237.2,
  230.4,
  224.8,
  223.4,
  223.9,
  224.2,
  226.6,
  229.1,
  229,
  228.2,
  220.3,
  227.7,
  232.6,
  232.7,
  233.8,
  232.8,
  231.9,
  231.6,
  326.4,
  273.1,
  237.8,
  234.2,
  232.7,
  230.8,
  228.5,
  227.5,
  227.4,
  226.6,
  225.5,
  225,
  224.6,
  223.8,
  222.5,
  221.2,
  220.9,
  220.9,
  219.9,
  218.4,
  218.2,
  218.8,
  219.2,
  219.7,
  219.8,
  219.1,
  221.1,
  223.1,
  222.8,
  221.6,
  223.2,
  221.2,
  218.2,
  219.1,
  222.2,
  222.9,
  225.6,
  229.4,
  229.3,
  229.6,
  221.5,
  229.6,
  233.6,
  234.5,
  234.9,
  234.9,
  234.7,
  234.3,
  324,
  270.9,
  237.8,
  234,
  232.1,
  231.7,
  232.3,
  233,
  232.7,
  230.6,
  230.4,
  228.9,
  228.2,
  226,
  225.4,
  224.7,
  225.2,
  228.7,
  230.2,
  226.8,
  228.2,
  231.9,
  226.4,
  226.7,
  231.1,
  241.5,
  237.2,
  239.5,
  241.6,
  237.1,
  238,
  240.1,
  230.3,
  229.6,
  238.7,
  245.5,
  242.1,
  235.3,
  235.8,
  236.1,
  232,
  243.2,
  259.5,
  261.2,
  256.8,
  258.4,
  254,
  260.1,
  285.8,
  261.2,
  270.7,
  291.8,
  298.4,
  285,
  287.9,
  275.1,
  245.9,
  242.1,
  240.4,
  236.8,
  238,
  239.4,
  240.7,
  243.2,
  268.9,
  302.5,
  269.5,
  252.3,
  254,
  260.5,
  300.1,
  287.6,
  265.4,
  263.6,
  290.6,
  311.6,
  311.1,
  310.7,
  306.6,
  302.5,
  303.8,
  308.5,
  308.3,
  305.9,
  309.1,
  314.2,
  316.2,
  316.7,
  303.2,
  296,
  307.6,
  319.5,
  325,
  328.2,
  321.8,
  307.7,
  350.4,
  305.1,
  267.5,
  267.5,
  266.5,
  265.3,
  264.6,
  262.6,
  263.3,
  262.6,
  264.7,
  262,
  260,
  260.2,
  259.4,
  259.1,
  259.5,
  257.5,
  257.1,
  256.4,
  256.2,
  257,
  255.5,
  256.3,
  257.6,
  251.1,
  250.6,
  252.8,
  255.1,
  255.6,
  254.9,
  254.2,
  250.3,
  249.8,
  250.5,
  252,
  253.3,
  255.7,
  256.8,
  258.5,
  253.7,
  261.2,
  266.4,
  267.5,
  267.2,
  266.5,
  265.4,
  264.2,
  339.4,
  290.6,
  263.2,
  261.1,
  259.6,
  259.7,
  259.5,
  258.4,
  257.6,
  257.7,
  258.9,
  254.1,
  253,
  252.9,
  251.9,
  250.2,
  251.7,
  257.9,
  288.8,
  317,
  321.2,
  321.3,
  321.4,
  322,
  321.7,
  321.9,
  322,
  322,
  322,
  321.7,
  322.6,
  322.1,
  320.9,
  321.5,
  321.8,
  321.7,
  321.9,
  322,
  322.2,
  322.7,
  321.9,
  322,
  316.8,
  293.9,
  270.5,
  252,
  251.2,
  249.9,
  322,
  277.6,
  249,
  250.7,
  252.4,
  251.4,
  250.8,
  252.5,
  254.1,
  251.9,
  251.2,
  252.9,
  252.5,
  257.4,
  266.7,
  289.2,
  288.4,
  300.1,
  306.2,
  307.5,
  308.3,
  308.9,
  312.3,
  312.7,
  312.9,
  313.4,
  313.3,
  313.3,
  313.8,
  313.9,
  313.5,
  313.2,
  313.4,
  314.7,
  314.4,
  314.2,
  316.3,
  318.5,
  319.8,
  322.6,
  323.3,
  325.5,
  327.2,
  331.4,
  333.8,
  334.7,
  336.4,
  337.2,
  351.7,
  343.4,
  340.5,
  340.8,
  339.3,
  337,
  336.6,
  336.5,
  335.9,
  334.3,
  334,
  334,
  334.9,
  335.4,
  335.4,
  334.2,
  336.2,
  335.5,
  333.9,
  329.3,
  332.4,
  333.3,
  333.5,
  332.8,
  332.3,
  331.5,
  331.2,
  330.5,
  328.7,
  330.6,
  330.1,
  330.8,
  330.9,
  330.8,
  330.2,
  330.3,
  332.3,
  333,
  333,
  334.3,
  332.2,
  341.1,
  346.7,
  345.5,
  344.3,
  342.1,
  340,
  335.2,
  355,
  340.5,
  331.5,
  324.4,
  310,
  295.1,
  287.8,
  264.2,
  258.3,
  257.2,
  255.8,
  254.2,
  252.1,
  251.2,
  251,
  250.3,
  250.3,
  250.1,
  249.6,
  248.8,
  247.8,
  247.4,
  247,
  246.7,
  245.8,
  245.6,
  245.5,
  245.6,
  244.7,
  244.2,
  243.4,
  242.2,
  238.1,
  236.8,
  236.8,
  238.3,
  240.8,
  242.3,
  244.4,
  246.1,
  243.3,
  249.9,
  256.4,
  258.9,
  259.1,
  259.3,
  263.1,
  263.5,
  310,
  269.8,
  261.8,
  263.7,
  292.3,
  293.8,
  309,
  288.6,
  308.1,
  333.1,
  341.7,
  340.2,
  346.3,
  347.2,
  347.7,
  347.7,
  343.5,
  340.2,
  340.5,
  341.3,
  341.9,
  342.8,
  344.4,
  345.3,
  346.7,
  348.1,
  348.8,
  350.3,
  352.2,
  353.5,
  355.3,
  356,
  358.1,
  359.5,
  362.4,
  368,
  370.4,
  371.6,
  375.7,
  379.3,
  363.2,
  325.3,
  333.5,
  362.1,
  358.9,
  347.6,
  343.3,
  367.4,
  380.6,
  334.3,
  333.3,
  308.9,
  304.6,
  296.7,
  295.7,
  298.9,
  301.7,
  303.5,
  308.7,
  308.1,
  310.7,
  323.4,
  328.8,
  337.6,
  339.5,
  330.5,
  332.4,
  335.5,
  341.8,
  360.2,
  353.5,
  354.6,
  356.5,
  359.9,
  361.9,
  364.7,
  364.5,
  362.3,
  360.9,
  363,
  364,
  367.6,
  369.6,
  370.6,
  373.4,
  376,
  376.9,
  377.7,
  378,
  378.1,
  377,
  365,
  359.1,
  359.3,
  364,
  353.8,
  343.3,
  300.1,
  327.3,
  295.8,
  298.3,
  294.7,
  310.1,
  335.9,
  337.8,
  341.3,
  346.6,
  351,
  362.2,
  363.8,
  366.5,
  368.4,
  369.6,
  369.1,
  368.7,
  367.9,
  365.5,
  366.3,
  366.4,
  361.4,
  350.4,
  365.1,
  368.9,
  370.9,
  371.6,
  371.1,
  363,
  360.2,
  357.8,
  359.3,
  359.4,
  358.7,
  360.8,
  361.3,
  363.1,
  363,
  362.2,
  362.4,
  361.9,
  361.6,
  362,
  362.9,
  362.5,
  362.1,
  368.4,
  363,
  361.9,
  361.5,
  361.6,
  357.8,
  354.4,
  349.9,
  343.1,
  298.3,
  280.1,
  315.7,
  301,
  323.3,
  303.2,
  277.7,
  276.2,
  291.1,
  315.9,
  329.1,
  312.8,
  299,
  332.1,
  296.6,
  277.7,
  277.1,
  281.6,
  295,
  307,
  281,
  290.3,
  283,
  310.1,
  316.8,
  338.6,
  350.8,
  352,
  348.5,
  324.2,
  350.7,
  342.9,
  333.1,
  357.3,
  357.6,
  344.5,
  316.4,
  305.6,
  290.5,
  338.3,
  290.8,
  284,
  296.2,
  334.6,
  315.8,
  280.5,
  275.7,
  273.1,
  273.1,
  282.3,
  283.1,
  292.4,
  310.3,
  340.5,
  344,
  351.2,
  350.5,
  351.9,
  360.1,
  359.1,
  359,
  359.1,
  359.8,
  360.1,
  360.4,
  360.7,
  361,
  360.7,
  359.5,
  358.7,
  354.8,
  352.7,
  350.8,
  354.6,
  361.6,
  346.2,
  279.2,
  287.1,
  292.9,
  285.9,
  314.6,
  324.2,
  319.9,
  323.1,
  316,
  303.7,
  275.3,
  295.5,
  291.3,
  274.3,
  274.1,
  272.5,
  271.1,
  269.9,
  269.5,
  277.8,
  274.7,
  268.1,
  269.8,
  279,
  270.9,
  293.6,
  340.9,
  340.4,
  345.2,
  345.9,
  343.9,
  338.4,
  300.6,
  268,
  265.3,
  265.6,
  266.8,
  270.9,
  267.2,
  272.5,
  324.3,
  343.8,
  344.1,
  343.3,
  342.3,
  344,
  345.5,
  346.5,
  347.2,
  345.7,
  341.4,
  348.6,
  316.5,
  315.7,
  312.1,
  310.9,
  317.8,
  313.4,
  339.6,
  341.1,
  334.7,
  337.8,
  352.2,
  355.8,
  355.4,
  355.3,
  355.6,
  355.7,
  355.8,
  355.1,
  353.6,
  352.6,
  353.1,
  351.8,
  349.3,
  351.1,
  351.8,
  351,
  350.9,
  352.1,
  351.5,
  350.7,
  350.8,
  349.3,
  343.7,
  325.5,
  292.4,
  274.6,
  260.3,
  260.1,
  260.2,
  284.1,
  330.5,
  338.4,
  338.8,
  339.6,
  342.6,
  344.2,
  342.7,
  344.6,
  345.8,
  346.8,
  348.7,
  348.8,
  347.7,
  346.9,
  345.8,
  350,
  351.1,
  345.2,
  345.4,
  346.3,
  346.7,
  346,
  346.3,
  345.9,
  343.6,
  343.2,
  345.5,
  347.4,
  349,
  349.5,
  347.4,
  344.6,
  342.9,
  341,
  339.1,
  338.9,
  338.8,
  340.9,
  338.7,
  336.6,
  336.4,
  336.4,
  336.4,
  334.8,
  332.2,
  332.4,
  337.5,
  333.8,
  333.4,
  330.1,
  330.3,
  337.5,
  342.1,
  344,
  356.2,
  359.5,
  360.6,
  362.6,
  364.1,
  363.4,
  362.1,
  359.9,
  390,
  368.6,
  356.1,
  348.9,
  346.9,
  346.4,
  344.8,
  342.5,
  339.5,
  337.4,
  337,
  337.6,
  338.3,
  338.4,
  339.4,
  339.3,
  338.4,
  338.4,
  339.3,
  340,
  340.1,
  340.2,
  340.5,
  341.4,
  341.1,
  340.1,
  339.4,
  338.2,
  337.8,
  337.1,
  337.1,
  336.5,
  336.5,
  337,
  337.1,
  337.8,
  339.6,
  341.2,
  341.9,
  341.9,
  343.8,
  344.6,
  345.4,
  345.6,
  345.6,
  344.4,
  341.6,
  335.2,
  356.1,
  341.4,
  338.4,
  338.1,
  337.1,
  337.7,
  337.6,
  338.1,
  338.5,
  339.5,
  339.8,
  338.8,
  337.9,
  335.7,
  333.8,
  326.4,
  334.4,
  334.7,
  331.6,
  326.4,
  261.8,
  310.8,
  331.7,
  331.2,
  330.4,
  326.3,
  328.4,
  287.8,
  274.7,
  298,
  266.5,
  277.2,
  291.5,
  308.7,
  318,
  286.8,
  268.1,
  263.6,
  262.5,
  275.7,
  289.5,
  337.8,
  341.8,
  342.4,
  343.5,
  344.2,
  344.7,
  343.5,
  352.9,
  346.6,
  342.9,
  340.9,
  340.9,
  339.2,
  319.7,
  299.8,
  279,
  325,
  277.3,
  297,
  333.3,
  341.4,
  338.9,
  337.4,
  331.3,
  329.5,
  328,
  346,
  347.8,
  348.4,
  348.7,
  347.3,
  346.3,
  348.6,
  349.9,
  349.2,
  349.4,
  349.5,
  350.5,
  351,
  351.4,
  352.4,
  353.1,
  353.8,
  355.1,
  355.9,
  357.1,
  357.9,
  358.8,
  359.5,
  360.3,
  360.9,
  361.6,
  363.1,
  363.4,
  363.7,
  370.4,
  365.8,
  364.3,
  364.1,
  364.4,
  365,
  365.7,
  365.7,
  365.7,
  366.2,
  366.3,
  366.2,
  366.7,
  366.7,
  366.9,
  367.4,
  367.4,
  367.5,
  368.7,
  369.8,
  369.6,
  367.9,
  367.8,
  367.8,
  367.6,
  367.5,
  367.5,
  367.4,
  367.2,
  367.7,
  367.3,
  367.3,
  367.2,
  366.8,
  367.6,
  368.5,
  369.2,
  370.2,
  371.5,
  373,
  372.6,
  372.3,
  370.7,
  368.1,
  364.8,
  363.9,
  363.2,
  360.7,
  383.2,
  355.9,
  348.9,
  353.2,
  341.4,
  330.6,
  308.6,
  296.1,
  278.6,
  278.5,
  278.7,
  280.2,
  280.2,
  284.5,
  284.7,
  272.5,
  271.6,
  274.1,
  277.1,
  272.2,
  267.8,
  271.1,
  274.4,
  276.1,
  276.3,
  277.6,
  278.2,
  277.1,
  274,
  271.8,
  269.2,
  265.4,
  260.9,
  255.7,
  249,
  245.8,
  245.9,
  246.6,
  247.2,
  246.8,
  248.3,
  244.3,
  251.3,
  255.9,
  257.5,
  257.5,
  256.3,
  256.1,
  304.6,
  267.4,
  253.5,
  253,
  253,
  256.2,
  257.5,
  255.7,
  254.6,
  252.9,
  251.3,
  250.2,
  247.7,
  246.4,
  244.7,
  242.3,
  240.4,
  239.7,
  241,
  241,
  241.2,
  240.5,
  240.4,
  239.9,
  239.8,
  240.3,
  240.4,
  240.5,
  240.8,
  241.2,
  241.9,
  241.6,
  241.9,
  241.8,
  240,
  239.7,
  241.5,
  244.1,
  246.5,
  247.6,
  248.1,
  243,
  248.2,
  253.6,
  254.9,
  254.8,
  255.5,
  256.3,
  298.6,
  271.2,
  255.4,
  254.8,
  253.3,
  250.9,
  249.4,
  247.3,
  247.2,
  247.2,
  246.8,
  246.7,
  247.7,
  251.4,
  256.1,
  262.4,
  265.4,
  267.3,
  265.1,
  261.5,
  261.5,
  262.2,
  261.2,
  265.2,
  314.4,
  299.2,
  260.9,
  251.2,
  248.1,
  243.8,
  240.6,
  239.5,
  240.7,
  246.8,
  236.4,
  233,
  233.6,
  234.4,
  234.4,
  234.2,
  233.7,
  226.8,
  231.8,
  236.5,
  237.6,
  237.3,
  236.8,
  236.5,
  294.4,
  246.2,
  235.8,
  233.6,
  232,
  230.4,
  229.8,
  228.1,
  226.4,
  225.5,
  225.4,
  226.5,
  227.2,
  228.1,
  231.5,
  295.9,
  307.5,
  318.2,
  281.6,
  268.5,
  282.8,
  286.8,
  290.9,
  305.4,
  319.6,
  320.8,
  319.7,
  320.6,
  323.1,
  323.5,
  324.3,
  324.4,
  319.1,
  316.3,
  313.8,
  313,
  314.3,
  316.2,
  318.9,
  317.7,
  320.4,
  324.4,
  316.9,
  300.3,
  318.1,
  328.2,
  329.5,
  331.2,
  338.7,
  338.8,
  332.8,
  331.2,
  331.2,
  318.2,
  292.1,
  315.1,
  329.4,
  328.5,
  328.7,
  332.7,
  332.2,
  335.5,
  339.2,
  333.7,
  318.9,
  337.3,
  318.6,
  314.5,
  331.9,
  331.5,
  330.1,
  344.6,
  345.1,
  347.3,
  347.5,
  348.2,
  345.1,
  331.5,
  327,
  346.4,
  347.1,
  347.6,
  343.8,
  340.9,
  331.7,
  334.2,
  340.3,
  348.3,
  351.1,
  353.7,
  353.3,
  351.4,
  350.7,
  354.1,
  354,
  354,
  362.1,
  360.1,
  352.7,
  353.3,
  354.1,
  343.8,
  332,
  342.8,
  351.6,
  345,
  343.7,
  347,
  349.3,
  350.1,
  349.4,
  349.2,
  349.9,
  350.2,
  349.5,
  347.8,
  349.7,
  349.6,
  349.2,
  348.1,
  345.5,
  347.7,
  346.4,
  344.8,
  343.5,
  342.2,
  342,
  343,
  342.7,
  342.6,
  341.2,
  339.8,
  336.8,
  339,
  343.1,
  339.8,
  340.2,
  345,
  345.4,
  344.4,
  344.6,
  342,
  333.9,
  300.5,
  329.1,
  302.6,
  303,
  291.8,
  286.4,
  328.4,
  339.4,
  341.2,
  341.3,
  341.7,
  341.8,
  342.4,
  342,
  342.3,
  340.7,
  338.5,
  325.6,
  306.1,
  300.2,
  313,
  332.2,
  333.1,
  332.1,
  313.2,
  304,
  303.9,
  322.1,
  320.7,
  319.7,
  331.9,
  334.6,
  335.2,
  334.5,
  333.8,
  334,
  333.5,
  334,
  333.8,
  333.7,
  334.6,
  334.9,
  335.6,
  335.1,
  336.3,
  337.7,
  338.4,
  339,
  338.7,
  351.8,
  340.9,
  337.5,
  336.8,
  336.5,
  335.8,
  334.8,
  334.7,
  334.9,
  335.2,
  335.4,
  334.8,
  333.7,
  334.7,
  335.7,
  336.2,
  335.8,
  336,
  335.8,
  335.3,
  334.9,
  334.9,
  334,
  333.6,
  331,
  329,
  326,
  323.8,
  324,
  324.3,
  324,
  323.2,
  322.5,
  320.8,
  319.1,
  319.1,
  318.8,
  319,
  319.9,
  320.5,
  320.3,
  318.2,
  309.8,
  304.8,
  299.1,
  305.3,
  312.7,
  316.1,
  327.6,
  305.1,
  269.4,
  264.8,
  279.5,
  279.8,
  275.9,
  266.7,
  260.2,
  252.5,
  261.4,
  273,
  283.4,
  292.2,
  269.6,
  272.4,
  263.9,
  259.5,
  265.1,
  255.6,
  252.2,
  247.3,
  252,
  247.3,
  243.3,
  243.1,
  244.6,
  252.5,
  268.1,
  279,
  283,
  289.3,
  291.9,
  296.6,
  272.3,
  249.6,
  251.1,
  265.4,
  270.2,
  266.7,
  263.6,
  267.5,
  268,
  270.6,
  273.6,
  268,
  260.9,
  261.7,
  295.3,
  319.7,
  304.9,
  270.8,
  264.7,
  267.5,
  268.2,
  268.9,
  272.5,
  305.3,
  303.7,
  286.3,
  301.6,
  303.2,
  301.9,
  273.9,
  262.7,
  261.7,
  261.7,
  261.4,
  260.3,
  260.1,
  260.4,
  288.1,
  317,
  304.2,
  301.9,
  264.4,
  258.8,
  258.3,
  257.8,
  256.9,
  258.3,
  258.3,
  262.5,
  280.7,
  300.8,
  313.4,
  314.5,
  315.9,
  316,
  314.7,
  314.5,
  319.7,
  309.5,
  310,
  316.4,
  324.3,
  340.8,
  326.9,
  323.4,
  322.3,
  310.3,
  322.7,
  326.1,
  324.6,
  325,
  325.3,
  321.1,
  321.9,
  316,
  315.7,
  317.3,
  318.6,
  317.3,
  322.3,
  323.2,
  322.1,
  324.1,
  327.4,
  329.2,
  326.6,
  327.7,
  325.8,
  326.2,
  327.2,
  325.6,
  319.6,
  319.6,
  324.5,
  326.3,
  324.5,
  327.6,
  329.2,
  329.1,
  328.1,
  330.1,
  324.2,
  328.1,
  329.8,
  328,
  332.9,
  335.6,
  335.8,
  336.7,
  336.4,
  341.7,
  337.9,
  334.7,
  335,
  333,
  334.2,
  336.9,
  336.2,
  337,
  337.5,
  338,
  337.6,
  337,
  336.6,
  335.9,
  335.7,
  336.1,
  336,
  335.6,
  335.5,
  335.3,
  335.4,
  335.7,
  335.9,
  336.3,
  336.5,
  337.1,
  337.3,
  337.8,
  337.7,
  338.4,
  338.3,
  338.9,
  339.8,
  340.3,
  341.5,
  342.3,
  343,
  343.3,
  344.3,
  344.8,
  342.9,
  339,
  339.2,
  340.6,
  344.2,
  346.6,
  344.9,
  351.1,
  346.4,
  345.4,
  347.4,
  348.5,
  349.1,
  350.1,
  351.3,
  352.2,
  353.4,
  354.7,
  351.4,
  354.1,
  352.1,
  353.7,
  351.5,
  321.5,
  325.4,
  331.7,
  322.5,
  340.9,
  351.2,
  354.7,
  352.4,
  352.7,
  352.3,
  353,
  355.6,
  357.7,
  358.3,
  357.7,
  357.7,
  356.6,
  356.2,
  357.7,
  356.7,
  358,
  353.9,
  355.3,
  359.3,
  359.3,
  356.9,
  360.5,
  359.9,
  358.1,
  349.7,
  360.7,
  356.1,
  349.4,
  326.5,
  353.4,
  351.2,
  351,
  348.6,
  345.8,
  351.5,
  349.4,
  348.2,
  347.3,
  342.8,
  331.8,
  340.9,
  305.3,
  291.7,
  298.3,
  294.7,
  316.5,
  313,
  326.6,
  334.9,
  336.2,
  336.9,
  337.3,
  340.3,
  333.2,
  332.8,
  343.4,
  345.2,
  346.3,
  347.9,
  349.6,
  349.9,
  350.4,
  351,
  350.6,
  349.8,
  347.6,
  351.9,
  354.8,
  354.7,
  354.3,
  354.8,
  353.9,
  353.2,
  353.3,
  352.3,
  355.9,
  351,
  351.1,
  351.9,
  347.2,
  347,
  345.4,
  346.7,
  348.5,
  344.5,
  341.3,
  339.6,
  338.5,
  337.5,
  338,
  337,
  337,
  336.2,
  335.5,
  322.9,
  320.8,
  319.2,
  317.1,
  315.9,
  314.8,
  312.2,
  310.3,
  308.3,
  304.8,
  302.3,
  298.4,
  295.7,
  288.4,
  267.3,
  247.9,
  242.7,
  247.6,
  244,
  239.6,
  242.8,
  245.8,
  240,
  246.9,
  253.8,
  260.9,
  271.4,
  260.7,
  279.2,
  338.7,
  273.6,
  260.8,
  292.8,
  269.3,
  254,
  269.3,
  294.5,
  255.4,
  259.4,
  285.1,
  276.4,
  291.5,
  312.7,
  318.7,
  319.7,
  319.4,
  321.2,
  324.2,
  327.5,
  326.6,
  326.1,
  325.7,
  325.3,
  326.3,
  327.7,
  326.1,
  323.7,
  321.9,
  320.7,
  319.4,
  318.5,
  318,
  317.9,
  317.4,
  317.6,
  317.2,
  318.3,
  319.2,
  320.8,
  308,
  290.6,
  286.7,
  285.6,
  283.1,
  281.4,
  280.7,
  282,
  296.3,
  283,
  282,
  281.4,
  281.5,
  279.9,
  273.2,
  272,
  272.3,
  272,
  268.6,
  269.1,
  270.9,
  272.6,
  274.9,
  296.4,
  305.3,
  311.9,
  311.6,
  313.4,
  311.7,
  311.2,
  305.7,
  284.6,
  276.7,
  266.3,
  264.4,
  264.6,
  257.3,
  253.6,
  247.9,
  239.7,
  238.1,
  236.5,
  236.7,
  233,
  233.9,
  234.2,
  238.1,
  242.9,
  246.8,
  239.3,
  248.9,
  257.3,
  285.9,
  307.6,
  282.9,
  265.8,
  303.3,
  310.3,
  303.8,
  307.4,
  306.2,
  307.2,
  300.6,
  304.1,
  308.1,
  308.2,
  309.2,
  310.5,
  312.7,
  310.2,
  312.3,
  307.3,
  306.1,
  302,
  269.3,
  243.8,
  244.5,
  242,
  257.3,
  295.3,
  313.9,
  313.9,
  314.5,
  314.2,
  315.6,
  315.3,
  315.7,
  316.9,
  317.9,
  318.6,
  310.9,
  287.3,
  283.1,
  288.2,
  303.4,
  312.4,
  313.9,
  316.8,
  316.7,
  315.5,
  313.6,
  314.8,
  313,
  312,
  318.7,
  300.7,
  244.5,
  238.1,
  236.3,
  233.2,
  232.7,
  234.1,
  236.6,
  233.8,
  235.2,
  237.5,
  237.9,
  238.7,
  239,
  244.1,
  267.3,
  270.4,
  251.2,
  282.6,
  249.8,
  248.1,
  272,
  281.3,
  299,
  298,
  298,
  294.6,
  297,
  295,
  288,
  271.2,
  268.9,
  301.2,
  277.3,
  283.5,
  304.4,
  318.2,
  320,
  322.9,
  324.6,
  325.7,
  324.1,
  319.5,
  317.6,
  295.9,
  280.9,
  291.5,
  313.5,
  310.7,
  298,
  294.1,
  300.5,
  302.2,
  257.8,
  254.8,
  246.9,
  247.2,
  247.4,
  248.9,
  249.8,
  250.2,
  248.5,
  244.5,
  244,
  244.1,
  247.7,
  247.7,
  247.8,
  249.7,
  249.5,
  249.2,
  253.3,
  266.6,
  291.2,
  314.3,
  311.8,
  294.5,
  314.4,
  302.3,
  300.6,
  306.4,
  308.8,
  310.9,
  322.3,
  323.8,
  320.9,
  321.7,
  324.8,
  324.7,
  324.5,
  325.3,
  327,
  326.8,
  327.4,
  328.2,
  330.6,
  330.2,
  330.3,
  331.4,
  331.8,
  333.7,
  335,
  336.3,
  337.7,
  338.1,
  339.3,
  339.5,
  339.8,
  340.3,
  340.2,
  340.2,
  340.7,
  340.1,
  339.9,
  339.5,
  337.2,
  337.9,
  337,
  328.5,
  312.6,
  306.5,
  287.6,
  317.2,
  324.9,
  326.1,
  327.6,
  328.3,
  327.4,
  324.8,
  318.6,
  297.8,
  286.5,
  315.1,
  318.9,
  319.5,
  320.7,
  321.8,
  322.9,
  323.8,
  322,
  276.9,
  266.5,
  266.3,
  278.6,
  261.3,
  255.2,
  254.1,
  256.1,
  253.1,
  261.1,
  258,
  256.6,
  250.3,
  252.5,
  257.5,
  263.1,
  266.9,
  272.7,
  280.4,
  272.1,
  253.5,
  236.5,
  236,
  242.6,
  293,
  285,
  321.8,
  339,
  340.7,
  341.1,
  341.5,
  339.8,
  337.4,
  332.2,
  332.9,
  335.3,
  335.2,
  333.5,
  335.1,
  334,
  334.1,
  335.7,
  336.4,
  337.5,
  337.2,
  337.2,
  337.6,
  338.2,
  338.8,
  339.3,
  339.9,
  346.5,
  345.2,
  344.5,
  345.4,
  346.8,
  324.7,
  302,
  299.7,
  344.6,
  339.8,
  348.4,
  350,
  348.3,
  334.8,
  348.6,
  351,
  351.5,
  351.5,
  351.7,
  353.5,
  353.2,
  344.7,
  328.5,
  349.1,
  334.4,
  329.5,
  336.7,
  348.1,
  353,
  353.2,
  337.4,
  327.6,
  344.2,
  345.4,
  326.2,
  335,
  345.6,
  349.5,
  343.7,
  333.5,
  320.7,
  287.1,
  305.4,
  336.5,
  335.6,
  336.5,
  340,
  314.3,
  324.1,
  319.4,
  330.9,
  315.6,
  339.6,
  347.5,
  351.9,
  355.7,
  356,
  354.9,
  355.4,
  356,
  357.4,
  357.9,
  359,
  362.4,
  363.6,
  363.4,
  362.9,
  363.5,
  362.5,
  363.5,
  365.4,
  365.9,
  367.1,
  367.8,
  367.9,
  367.6,
  367.9,
  366.9,
  365.1,
  363.2,
  362.4,
  361.8,
  362.4,
  360.4,
  348.7,
  359.5,
  363.9,
  364.4,
  363.7,
  364.8,
  364.9,
  366.7,
  368.4,
  369.2,
  370.7,
  372.3,
  377.7,
  374.8,
  370.7,
  365.1,
  367,
  324,
  302.3,
  310.6,
  336,
  354.3,
  357.9,
  361.9,
  360.9,
  359.5,
  355.6,
  352.3,
  353.3,
  338.6,
  351.1,
  340.7,
  343.5,
  320.8,
  325.1,
  351.6,
  331.1,
  324.8,
  349.4,
  346.7,
  354.8,
  367.9,
  367.4,
  367.1,
  366.9,
  364.7,
  368.2,
  368,
  368.4,
  368.2,
  368.7,
  369.3,
  369.4,
  373.2,
  356.7,
  368.9,
  365.3,
  332.5,
  344.5,
  330.6,
  368.2,
  356.7,
  354.9,
  345.7,
  336.3,
  342.9,
  340.8,
  356.2,
  359.8,
  347.4,
  364.7,
  363.5,
  356.7,
  363.2,
  361.7,
  350.3,
  348.7,
  339.2,
  326.7,
  349.6,
  350.9,
  354.8,
  355,
  356.4,
  356,
  351.8,
  347,
  347.2,
  341.5,
  348.2,
  354.3,
  354.4,
  352.2,
  352.7,
  351.2,
  346.7,
  346.6,
  344.8,
  342.8,
  343.7,
  345,
  346.2,
  348.5,
  343.8,
  340.8,
  342,
  338.8,
  330.2,
  350.9,
  347.8,
  342.5,
  324.8,
  344.3,
  347.3,
  344.8,
  341.1,
  336.8,
  334.5,
  337.2,
  320,
  305.3,
  300.3,
  303.9,
  330.2,
  302,
  277.6,
  257.8,
  264.8,
  264.9,
  262.5,
  254.3,
  251.7,
  281.3,
  295.2,
  274,
  292.9,
  301.7,
  318.3,
  323,
  284,
  261.6,
  276,
  287,
  292,
  282.7,
  282.8,
  259.2,
  256.9,
  259.2,
  264.7,
  290.4,
  315.8,
  322,
  330.9,
  345.4,
  351.6,
  363.4,
  355.7,
  351.6,
  351.4,
  350.9,
  351.4,
  350.2,
  348,
  349.7,
  349.3,
  346.4,
  340.9,
  331.9,
  337.1,
  338.6,
  341.1,
  338.9,
  339.8,
  339.5,
  338.7,
  340.4,
  337.4,
  338.7,
  337.3,
  337.6,
  336.4,
  335.3,
  336.6,
  335.1,
  334.1,
  333.3,
  329.5,
  328.6,
  330.5,
  331.1,
  327.9,
  332.2,
  336.3,
  335.8,
  345.5,
  349.4,
  350.9,
  321.4,
  265.7,
  310.4,
  311.3,
  302.3,
  292.1,
  341.6,
  328,
  325.1,
  328.5,
  308.6,
  318.8,
  316,
  317.1,
  315.8,
  315.5,
  307.4,
  305.8,
  273.5,
  244.2,
  239.5,
  238,
  237.9,
  261.6,
  302.3,
  313.5,
  284.4,
  237.2,
  236.3,
  247.8,
  273.6,
  313.7,
  315.4,
  316.4,
  317.7,
  313.3,
  309.6,
  309,
  282.5,
  274.2,
  270.4,
  306.4,
  308.2,
  309.4,
  307.6,
  308.3,
  308.3,
  307.5,
  305.9,
  302.9,
  304.4,
  298.3,
  280.6,
  289.9,
  318.4,
  284,
  277.8,
  296.1,
  274.6,
  273.7,
  286.3,
  272.2,
  278.3,
  239.6,
  242.5,
  244.2,
  253.1,
  227,
  233.2,
  221.2,
  217.1,
  219.8,
  218.1,
  251.3,
  269.7,
  289.6,
  287.7,
  291.1,
  291.9,
  292.9,
  293.6,
  294.2,
  294.4,
  294.4,
  292.3,
  292,
  291.8,
  290.1,
  268.7,
  254.6,
  276.1,
  257.9,
  244.6,
  221.6,
  224.7,
  223.4,
  205,
  209.1,
  209.7,
  209.2,
  210,
  210.8,
  244.2,
  220,
  212.4,
  212,
  212.5,
  212.1,
  211.6,
  211.6,
  211.4,
  211.8,
  211.9,
  211.8,
  212.4,
  212.7,
  212.1,
  212.2,
  212,
  211.9,
  211.1,
  210.8,
  210,
  209.1,
  209.4,
  209.8,
  210.4,
  209.9,
  209.5,
  209.1,
  208.1,
  208.1,
  207.6,
  207.8,
  207.5,
  206.6,
  205.9,
  203.5,
  202.4,
  199.8,
  201,
  201.3,
  204.5,
  210.4,
  221.9,
  259.2,
  285.1,
  301.7,
  304.5,
  302.9,
  315.8,
  308.6,
  309.7,
  310.4,
  300.9,
  309.7,
  307.5,
  302,
  304.6,
  295.4,
  297.9,
  298.6,
  301.7,
  297.5,
  303.4,
  307.4,
  314.1,
  317,
  319.3,
  322.1,
  323.1,
  324.2,
  322.2,
  302.1,
  299.1,
  275.8,
  261.6,
  261.3,
  323.7,
  324.3,
  271.3,
  270.2,
  273,
  276.8,
  278.1,
  278.8,
  307.6,
  315.8,
  309.5,
  292.4,
  324.5,
  336,
  338.2,
  345.7,
  345.6,
  343.4,
  344.8,
  345.6,
  347.1,
  341.8,
  337.7,
  337.4,
  336.5,
  333.8,
  334.7,
  335.2,
  328.5,
  337.1,
  341.1,
  340.8,
  335.8,
  331,
  334,
  331.3,
  331.4,
  338.6,
  339.5,
  341.6,
  342,
  342.3,
  341.8,
  338.9,
  337.9,
  337.2,
  337.3,
  337.5,
  336.7,
  337.3,
  339,
  340,
  340.9,
  340.3,
  341.4,
  343.7,
  344.3,
  341.9,
  341.5,
  343.4,
  345.5,
  344.6,
  336.2,
  319.3,
  333.4,
  348.8,
  346.2,
  338.6,
  355.8,
  354.6,
  354.3,
  352.1,
  347.5,
  343.4,
  323.8,
  300,
  293.3,
  314.9,
  344,
  341,
  336.7,
  339.7,
  337.1,
  318.8,
  326.5,
  330.5,
  330.9,
  337.4,
  331,
  308.7,
  277.8,
  263.8,
  267.8,
  279.8,
  291.3,
  297.7,
  300.4,
  302.6,
  304.3,
  306.7,
  309.8,
  310.9,
  308.7,
  306.3,
  303.6,
  303.8,
  307.3,
  308,
  307.9,
  302.3,
  289.6,
  273.6,
  272.8,
  272.7,
  274.2,
  278,
  309.5,
  293.7,
  287.7,
  280.4,
  278.6,
  277.1,
  286.9,
  301.5,
  304.5,
  302.8,
  308,
  308,
  308.9,
  310.5,
  318.9,
  326.5,
  326.7,
  328.3,
  326.8,
  327.3,
  329.4,
  329.1,
  328.2,
  327.5,
  326.9,
  326.6,
  326.5,
  325.8,
  325.2,
  324.7,
  324.3,
  323.7,
  323.8,
  324.1,
  324,
  324.7,
  326.4,
  327.4,
  328.5,
  329.9,
  330.1,
  330.6,
  330.6,
  330.5,
  330.6,
  330.2,
  330.3,
  330,
  334.5,
  330.6,
  329.8,
  329.7,
  329.7,
  329.2,
  328.2,
  328.2,
  328.1,
  328,
  328,
  328.6,
  328.5,
  328.9,
  329.1,
  329,
  329.4,
  329.3,
  329.4,
  329.6,
  329.1,
  328.9,
  328.5,
  328.5,
  328.1,
  327.9,
  326.9,
  326.4,
  325.3,
  324.7,
  324.3,
  323.6,
  323.4,
  323.3,
  322.8,
  323.2,
  323.6,
  324.6,
  325.9,
  327.4,
  327.6,
  328.4,
  328.4,
  328.3,
  328,
  327,
  324.6,
  323.7,
  329.8,
  324.7,
  322.5,
  322.4,
  322.9,
  322,
  321.9,
  322.7,
  322.4,
  322.9,
  323.1,
  322.6,
  322.7,
  323,
  323.1,
  323.7,
  323,
  321.3,
  321.7,
  321.7,
  318.8,
  316,
  315.9,
  316.5,
  316.3,
  316.2,
  316,
  316.1,
  316.1,
  316.5,
  318.1,
  318.7,
  319.2,
  319.5,
  320.3,
  321,
  320.6,
  320.9,
  322.9,
  321.3,
  325.9,
  331,
  331.7,
  332,
  332.5,
  332.4,
  332.5,
  332.1,
  337.3,
  331.7,
  330.5,
  330.9,
  331.5,
  332.6,
  333.9,
  335.9,
  337,
  338.4,
  339.5,
  340.3,
  340.8,
  341.4,
  341.9,
  342.5,
  342.9,
  343.7,
  343.8,
  344.2,
  344.4,
  345.3,
  346,
  346.7,
  347.4,
  348.9,
  350.1,
  351.7,
  354.3,
  357.3,
  360.2,
  361.7,
  363.6,
  364.7,
  366.6,
  367.8,
  368.9,
  369.2,
  369.4,
  370,
  370.4,
  370.8,
  372.2,
  373,
  373.3,
  373.6,
  373.2,
  373.6,
  377,
  376.4,
  374.4,
  372.5,
  371.2,
  370.6,
  371.9,
  370.7,
  369.5,
  368.7,
  368.5,
  368.6,
  367.7,
  364.5,
  359.3,
  359.5,
  350,
  325,
  305.5,
  320.2,
  318.1,
  304.6,
  291,
  291.7,
  280.7,
  271.8,
  282.5,
  273.1,
  272.3,
  277.5,
  282,
  288.1,
  289.3,
  316.7,
  332,
  319,
  305.8,
  291.9,
  292.6,
  299.5,
  306.2,
  313.7,
  322.6,
  355.5,
  357.4,
  358.6,
  364,
  367.3,
  370.8,
  362.2,
  365.4,
  368.3,
  366.9,
  350.1,
  312.4,
  323.5,
  328.8,
  289.2,
  313.6,
  315.4,
  331.3,
  314.2,
  290.1,
  319.3,
  311.6,
  325,
  320.8,
  307.7,
  307.7,
  318.1,
  345.5,
  340.2,
  339.1,
  340.5,
  345.3,
  343.4,
  346.6,
  341.3,
  339.1,
  341.9,
  341.8,
  342.3,
  346.2,
  342,
  337.6,
  344.9,
  348.2,
  348,
  346.7,
  345.1,
  345.4,
  347.1,
  348,
  345.1,
  347.8,
  342.2,
  348.8,
  309.9,
  288.7,
  274.5,
  303.8,
  338.2,
  345.4,
  345.8,
  345,
  344.7,
  344.1,
  344.3,
  344,
  341.4,
  341.2,
  339.9,
  339.8,
  338.9,
  338.4,
  338.9,
  340.6,
  341.2,
  339.8,
  337.9,
  337.6,
  338.5,
  338.8,
  339.9,
  340.5,
  337.9,
  336.5,
  337.4,
  337.4,
  337,
  336.1,
  336.1,
  336.6,
  340.3,
  344.5,
  346.7,
  347.3,
  346.8,
  347.5,
  348.9,
  349.7,
  348.3,
  328.2,
  338.7,
  350.1,
  345.7,
  343.7,
  344.3,
  344.1,
  345.1,
  345.5,
  345.5,
  344.5,
  344.3,
  344.9,
  345.3,
  343.9,
  342.5,
  342.2,
  341.8,
  342.3,
  342.3,
  342.1,
  341.6,
  341.5,
  342.4,
  341.6,
  340.1,
  339.2,
  338.2,
  336,
  335.6,
  335.2,
  333.8,
  331.7,
  331.5,
  330.5,
  330,
  327.7,
  324.3,
  319.9,
  330.4,
  336.9,
  339.7,
  340.8,
  343.5,
  308,
  304.8,
  316.2,
  288.5,
  276.6,
  309.8,
  330.2,
  331.7,
  332.2,
  314.5,
  323.8,
  334.6,
  333.5,
  336.9,
  335.4,
  336,
  334.6,
  333.3,
  335,
  336.2,
  335.5,
  336.6,
  336.7,
  332.1,
  314.3,
  301.1,
  322.4,
  334.3,
  338.6,
  323.1,
  318.1,
  303.7,
  296.3,
  323.2,
  333.5,
  336.5,
  336.2,
  333.4,
  330.4,
  328.3,
  326,
  325.8,
  328.9,
  333.6,
  337.6,
  323,
  265.3,
  244.3,
  240.6,
  250.9,
  255.1,
  262.2,
  273.8,
  308.1,
  322.3,
  335.3,
  337.6,
  340,
  341.9,
  342.4,
  342.7,
  343,
  343,
  340.6,
  341.1,
  339.9,
  338.4,
  337.3,
  337,
  336,
  335.1,
  335.3,
  333.8,
  331.5,
  331.2,
  330,
  330.6,
  329.8,
  328.3,
  327.4,
  325.7,
  309.6,
  282.7,
  264.5,
  281.5,
  287.3,
  303.5,
  312.1,
  305.4,
  316.3,
  323.5,
  318.8,
  297.5,
  285,
  311.9,
  325.7,
  327,
  294,
  306.7,
  299,
  284.6,
  331.2,
  357,
  348,
  344.7,
  344.8,
  348.5,
  348,
  341.1,
  344.7,
  344.7,
  349.5,
  349.3,
  346.3,
  346.4,
  344.5,
  340.5,
  340.2,
  344.8,
  345.7,
  345.6,
  344.4,
  340,
  337.3,
  347.9,
  336.5,
  343.2,
  347.3,
  332.4,
  296.4,
  328.8,
  346.8,
  347.4,
  352,
  353.2,
  353,
  354,
  354.1,
  354.4,
  355.9,
  357.4,
  357.3,
  358.4,
  358.8,
  358.6,
  357.8,
  356.3,
  351.3,
  344,
  344.5,
  359.6,
  341,
  346,
  338.7,
  324.6,
  322.4,
  334.3,
  332.3,
  320.6,
  326.1,
  327.7,
  325.2,
  315,
  307.8,
  307.4,
  313.8,
  312.3 ;

 CO2air =
  400,    400,   400,   400, 
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,    400,   400,   400,
  400,  400,  400,  400 ;

 hc =
  15.5 ;

 za =
  27 ;
}
