netcdf isnow_flg3l {
dimensions:
	x = 1;
	y = 1;
	tile = 17 ;
   msn = 3;
   ms = 6;
variables:
	integer isnow_flg3l(tile, y, x) ;
	float snow_rho1l(tile, y, x) ;
	float snage_tile(tile, y, x) ;
	float snow_rho1(tile, y, x) ;
	float snow_rho2(tile, y, x) ;
	float snow_rho3(tile, y, x) ;
	float snow_mass1(tile, y, x) ;
	float snow_mass2(tile, y, x) ;
	float snow_mass3(tile, y, x) ;
	float snow_depth1(tile, y, x) ;
	float snow_depth2(tile, y, x) ;
	float snow_depth3(tile, y, x) ;
	float snow_tmp1(tile, y, x) ;
	float snow_tmp2(tile, y, x) ;
	float snow_tmp3(tile, y, x) ;
	float sthu_tile1(tile, y, x) ;
	float sthu_tile2(tile, y, x) ;
	float sthu_tile3(tile, y, x) ;
	float sthu_tile4(tile, y, x) ;
	float sthu_tile5(tile, y, x) ;
	float sthu_tile6(tile, y, x) ;
	float sthf_tile1(tile, y, x) ;
	float sthf_tile2(tile, y, x) ;
	float sthf_tile3(tile, y, x) ;
	float sthf_tile4(tile, y, x) ;
	float sthf_tile5(tile, y, x) ;
	float sthf_tile6(tile, y, x) ;
	float smcl_tile1(tile, y, x) ;
	float smcl_tile2(tile, y, x) ;
	float smcl_tile3(tile, y, x) ;
	float smcl_tile4(tile, y, x) ;
	float smcl_tile5(tile, y, x) ;
	float smcl_tile6(tile, y, x) ;
	float tsoil_tile1(tile, y, x) ;
	float tsoil_tile2(tile, y, x) ;
	float tsoil_tile3(tile, y, x) ;
	float tsoil_tile4(tile, y, x) ;
	float tsoil_tile5(tile, y, x) ;
	float tsoil_tile6(tile, y, x) ;
data:

isnow_flg3l = 
0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ,  0, 0 ,  0, 0 , 0 , 0 , 0 ;

snow_rho1l = 
120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0;

snage_tile = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

snow_rho1 = 
120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0;

snow_rho2 = 
120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0;

snow_rho3 = 
120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0, 120.0;

snow_mass1 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

snow_mass2 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

snow_mass3 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

snow_depth1 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

snow_depth2 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

snow_depth3 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

snow_tmp1 = 
273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16;

snow_tmp2 = 
273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16;

snow_tmp3 = 
273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16,273.16;

sthu_tile1 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthu_tile2 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthu_tile3 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthu_tile4 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthu_tile5 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthu_tile6 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthf_tile1 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthf_tile2 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthf_tile3 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthf_tile4 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthf_tile5 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

sthf_tile6 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

smcl_tile1 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

smcl_tile2 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

smcl_tile3 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

smcl_tile4 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

smcl_tile5 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

smcl_tile6 = 
0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0;

tsoil_tile1 = 
280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0;

tsoil_tile2 = 
280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0;

tsoil_tile3 = 
280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0;

tsoil_tile4 = 
280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0;

tsoil_tile5 = 
280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0;

tsoil_tile6 = 
280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0, 280.0;

}
